
library ieee;
use ieee.std_logic_1164.all;
library work;
use work.cam_pkg.all;

entity romdata is
  generic (ADR_BITS  : integer;
           DATA_BITS : integer);             -- for compatibility
  port (
    clk : in  std_logic;
    a   : in  std_logic_vector(ADR_BITS-1 downto 0);
    q   : out std_logic_vector(DATA_BITS-1 downto 0));
end romdata;

architecture rtl of romdata is
    ATTRIBUTE ram_extract: string;
    ATTRIBUTE ram_extract OF q: SIGNAL IS "yes";
    ATTRIBUTE ram_style: string;
    ATTRIBUTE ram_style OF q: SIGNAL IS "block";
  
  signal areg : std_logic_vector((GRIDX_BITS+GRIDY_BITS-1) downto 0);  -- GRIDX+GRIDY-1
begin

  process(clk)
  begin
    if rising_edge(clk) then
      areg <= a(areg'high downto areg'low);
    end if;
  end process;

  process(areg)
  begin
    case areg is
      -- GRIDY+GRIDX --    REFY+REFX

when "000000000000" => q <= "00000000000000000000";
when "000000000001" => q <= "00000000000000001100";
when "000000000010" => q <= "00001010010010000001";
when "000000000011" => q <= "00011001010011010101";
when "000000000100" => q <= "00100100110100010001";
when "000000000101" => q <= "00101101100100111010";
when "000000000110" => q <= "00110100000101010100";
when "000000000111" => q <= "00111000110101100100";
when "000000001000" => q <= "00111100100101101100";
when "000000001001" => q <= "00111111000101101111";
when "000000001010" => q <= "01000000110101101111";
when "000000001011" => q <= "01000001110101101100";
when "000000001100" => q <= "01000010110101101000";
when "000000001101" => q <= "01000011010101100011";
when "000000001110" => q <= "01000011110101011110";
when "000000001111" => q <= "01000100000101011000";
when "000000010000" => q <= "01000100010101010011";
when "000000010001" => q <= "01000100110101001101";
when "000000010010" => q <= "01000101000101001000";
when "000000010011" => q <= "01000101100101000010";
when "000000010100" => q <= "01000110000100111101";
when "000000010101" => q <= "01000110100100110111";
when "000000010110" => q <= "01000111010100110010";
when "000000010111" => q <= "01001000000100101100";
when "000000011000" => q <= "01001000110100100110";
when "000000011001" => q <= "01001001100100100000";
when "000000011010" => q <= "01001010010100011001";
when "000000011011" => q <= "01001011000100010010";
when "000000011100" => q <= "01001011110100001100";
when "000000011101" => q <= "01001100100100000101";
when "000000011110" => q <= "01001100110011111111";
when "000000011111" => q <= "01001100110011111010";
when "000000100000" => q <= "01001100010011110110";
when "000000100001" => q <= "01001011000011110111";
when "000000100010" => q <= "01001000100011111100";
when "000000100011" => q <= "01000100100100001000";
when "000000100100" => q <= "00111110110100011111";
when "000000100101" => q <= "00110110110101000011";
when "000000100110" => q <= "00101011100101111100";
when "000000100111" => q <= "00011100100111000000";
when "000001000000" => q <= "00000000000000000000";
when "000001000001" => q <= "00000111110001011001";
when "000001000010" => q <= "00010111000010111100";
when "000001000011" => q <= "00100011000100000010";
when "000001000100" => q <= "00101100000100110010";
when "000001000101" => q <= "00110010100101010001";
when "000001000110" => q <= "00110111100101100100";
when "000001000111" => q <= "00111011000101101111";
when "000001001000" => q <= "00111101100101110011";
when "000001001001" => q <= "00111111000101110011";
when "000001001010" => q <= "01000000010101110000";
when "000001001011" => q <= "01000000110101101100";
when "000001001100" => q <= "01000001010101100110";
when "000001001101" => q <= "01000001100101100001";
when "000001001110" => q <= "01000001110101011011";
when "000001001111" => q <= "01000010000101010101";
when "000001010000" => q <= "01000010010101010000";
when "000001010001" => q <= "01000010100101001010";
when "000001010010" => q <= "01000010110101000101";
when "000001010011" => q <= "01000011010101000000";
when "000001010100" => q <= "01000011110100111011";
when "000001010101" => q <= "01000100010100110110";
when "000001010110" => q <= "01000100110100110001";
when "000001010111" => q <= "01000101100100101011";
when "000001011000" => q <= "01000110010100100101";
when "000001011001" => q <= "01000111010100011111";
when "000001011010" => q <= "01001000000100011001";
when "000001011011" => q <= "01001001000100010010";
when "000001011100" => q <= "01001010000100001011";
when "000001011101" => q <= "01001010110100000100";
when "000001011110" => q <= "01001011100011111100";
when "000001011111" => q <= "01001100000011110110";
when "000001100000" => q <= "01001100000011110000";
when "000001100001" => q <= "01001011100011101101";
when "000001100010" => q <= "01001010010011101110";
when "000001100011" => q <= "01000111110011110101";
when "000001100100" => q <= "01000011110100000100";
when "000001100101" => q <= "00111110000100100000";
when "000001100110" => q <= "00110101100101001100";
when "000001100111" => q <= "00101001110110001111";
when "000010000000" => q <= "00000100000000100000";
when "000010000001" => q <= "00010100000010010110";
when "000010000010" => q <= "00100000010011101011";
when "000010000011" => q <= "00101001110100100100";
when "000010000100" => q <= "00110000100101001011";
when "000010000101" => q <= "00110101110101100010";
when "000010000110" => q <= "00111001010101101111";
when "000010000111" => q <= "00111011110101110101";
when "000010001000" => q <= "00111101010101110110";
when "000010001001" => q <= "00111110100101110011";
when "000010001010" => q <= "00111111000101101111";
when "000010001011" => q <= "00111111100101101001";
when "000010001100" => q <= "00111111100101100100";
when "000010001101" => q <= "00111111110101011110";
when "000010001110" => q <= "00111111110101011000";
when "000010001111" => q <= "01000000000101010010";
when "000010010000" => q <= "01000000010101001101";
when "000010010001" => q <= "01000000010101001000";
when "000010010010" => q <= "01000000110101000011";
when "000010010011" => q <= "01000001000100111110";
when "000010010100" => q <= "01000001100100111001";
when "000010010101" => q <= "01000010000100110100";
when "000010010110" => q <= "01000010110100101111";
when "000010010111" => q <= "01000011010100101010";
when "000010011000" => q <= "01000100010100100101";
when "000010011001" => q <= "01000101000100011111";
when "000010011010" => q <= "01000110000100011001";
when "000010011011" => q <= "01000110110100010010";
when "000010011100" => q <= "01000111110100001011";
when "000010011101" => q <= "01001000110100000011";
when "000010011110" => q <= "01001001110011111011";
when "000010011111" => q <= "01001010100011110100";
when "000010100000" => q <= "01001011000011101101";
when "000010100001" => q <= "01001011010011101000";
when "000010100010" => q <= "01001010110011100101";
when "000010100011" => q <= "01001001010011100111";
when "000010100100" => q <= "01000110110011110001";
when "000010100101" => q <= "01000010100100000100";
when "000010100110" => q <= "00111100010100100111";
when "000010100111" => q <= "00110011010101011101";
when "000011000000" => q <= "00010000000001100001";
when "000011000001" => q <= "00011101000011001000";
when "000011000010" => q <= "00100110110100001111";
when "000011000011" => q <= "00101110010100111111";
when "000011000100" => q <= "00110011100101011101";
when "000011000101" => q <= "00110111010101101110";
when "000011000110" => q <= "00111001110101110110";
when "000011000111" => q <= "00111011100101111000";
when "000011001000" => q <= "00111100110101110110";
when "000011001001" => q <= "00111101010101110010";
when "000011001010" => q <= "00111101100101101101";
when "000011001011" => q <= "00111101110101100111";
when "000011001100" => q <= "00111101110101100000";
when "000011001101" => q <= "00111101110101011010";
when "000011001110" => q <= "00111110000101010101";
when "000011001111" => q <= "00111110000101001111";
when "000011010000" => q <= "00111110010101001010";
when "000011010001" => q <= "00111110100101000101";
when "000011010010" => q <= "00111110110101000000";
when "000011010011" => q <= "00111111000100111100";
when "000011010100" => q <= "00111111100100110111";
when "000011010101" => q <= "01000000000100110011";
when "000011010110" => q <= "01000000110100101110";
when "000011010111" => q <= "01000001010100101001";
when "000011011000" => q <= "01000010000100100100";
when "000011011001" => q <= "01000011000100011110";
when "000011011010" => q <= "01000011110100011000";
when "000011011011" => q <= "01000100110100010010";
when "000011011100" => q <= "01000101110100001011";
when "000011011101" => q <= "01000110110100000011";
when "000011011110" => q <= "01000111110011111011";
when "000011011111" => q <= "01001000110011110011";
when "000011100000" => q <= "01001001100011101011";
when "000011100001" => q <= "01001010000011100100";
when "000011100010" => q <= "01001010010011011111";
when "000011100011" => q <= "01001001100011011110";
when "000011100100" => q <= "01001000000011100010";
when "000011100101" => q <= "01000101010011110000";
when "000011100110" => q <= "01000000100100001010";
when "000011100111" => q <= "00111001110100110110";
when "000100000000" => q <= "00011000110010010101";
when "000100000001" => q <= "00100011010011101110";
when "000100000010" => q <= "00101011010100101011";
when "000100000011" => q <= "00110001000101010010";
when "000100000100" => q <= "00110101000101101001";
when "000100000101" => q <= "00110111110101110101";
when "000100000110" => q <= "00111001110101111010";
when "000100000111" => q <= "00111010110101111001";
when "000100001000" => q <= "00111011100101110110";
when "000100001001" => q <= "00111011110101110000";
when "000100001010" => q <= "00111100000101101010";
when "000100001011" => q <= "00111100000101100011";
when "000100001100" => q <= "00111100000101011101";
when "000100001101" => q <= "00111100000101010111";
when "000100001110" => q <= "00111100000101010001";
when "000100001111" => q <= "00111100010101001100";
when "000100010000" => q <= "00111100100101000111";
when "000100010001" => q <= "00111100110101000011";
when "000100010010" => q <= "00111101000100111110";
when "000100010011" => q <= "00111101100100111010";
when "000100010100" => q <= "00111101110100110110";
when "000100010101" => q <= "00111110010100110001";
when "000100010110" => q <= "00111111000100101101";
when "000100010111" => q <= "00111111100100101000";
when "000100011000" => q <= "01000000010100100011";
when "000100011001" => q <= "01000001000100011110";
when "000100011010" => q <= "01000001110100011000";
when "000100011011" => q <= "01000010110100010010";
when "000100011100" => q <= "01000011110100001011";
when "000100011101" => q <= "01000100110100000100";
when "000100011110" => q <= "01000101110011111100";
when "000100011111" => q <= "01000110110011110011";
when "000100100000" => q <= "01000111110011101010";
when "000100100001" => q <= "01001000100011100010";
when "000100100010" => q <= "01001001000011011011";
when "000100100011" => q <= "01001001000011010111";
when "000100100100" => q <= "01001000010011011000";
when "000100100101" => q <= "01000110010011100000";
when "000100100110" => q <= "01000011000011110011";
when "000100100111" => q <= "00111110000100010110";
when "000101000000" => q <= "00011111010010111111";
when "000101000001" => q <= "00100111110100001101";
when "000101000010" => q <= "00101110000101000000";
when "000101000011" => q <= "00110010100101100000";
when "000101000100" => q <= "00110101100101110010";
when "000101000101" => q <= "00110111110101111010";
when "000101000110" => q <= "00111001000101111011";
when "000101000111" => q <= "00111001110101111001";
when "000101001000" => q <= "00111010000101110100";
when "000101001001" => q <= "00111010010101101101";
when "000101001010" => q <= "00111010010101100110";
when "000101001011" => q <= "00111010010101100000";
when "000101001100" => q <= "00111010010101011001";
when "000101001101" => q <= "00111010010101010011";
when "000101001110" => q <= "00111010100101001110";
when "000101001111" => q <= "00111010110101001001";
when "000101010000" => q <= "00111010110101000101";
when "000101010001" => q <= "00111011010101000000";
when "000101010010" => q <= "00111011100100111100";
when "000101010011" => q <= "00111100000100111000";
when "000101010100" => q <= "00111100100100110100";
when "000101010101" => q <= "00111101000100110000";
when "000101010110" => q <= "00111101100100101100";
when "000101010111" => q <= "00111110000100100111";
when "000101011000" => q <= "00111110110100100010";
when "000101011001" => q <= "00111111010100011101";
when "000101011010" => q <= "01000000000100011000";
when "000101011011" => q <= "01000001000100010010";
when "000101011100" => q <= "01000001110100001011";
when "000101011101" => q <= "01000010110100000100";
when "000101011110" => q <= "01000011110011111100";
when "000101011111" => q <= "01000101000011110011";
when "000101100000" => q <= "01000110000011101010";
when "000101100001" => q <= "01000110110011100001";
when "000101100010" => q <= "01000111100011011001";
when "000101100011" => q <= "01000111110011010011";
when "000101100100" => q <= "01000111100011010001";
when "000101100101" => q <= "01000110100011010101";
when "000101100110" => q <= "01000100010011100010";
when "000101100111" => q <= "01000000100011111110";
when "000110000000" => q <= "00100100000011100001";
when "000110000001" => q <= "00101010110100100101";
when "000110000010" => q <= "00101111110101010000";
when "000110000011" => q <= "00110011010101101010";
when "000110000100" => q <= "00110101100101111000";
when "000110000101" => q <= "00110111000101111100";
when "000110000110" => q <= "00111000000101111011";
when "000110000111" => q <= "00111000100101110111";
when "000110001000" => q <= "00111000110101110001";
when "000110001001" => q <= "00111000110101101010";
when "000110001010" => q <= "00111000110101100011";
when "000110001011" => q <= "00111000110101011100";
when "000110001100" => q <= "00111000110101010110";
when "000110001101" => q <= "00111001000101010000";
when "000110001110" => q <= "00111001000101001011";
when "000110001111" => q <= "00111001010101000111";
when "000110010000" => q <= "00111001100101000010";
when "000110010001" => q <= "00111001110100111110";
when "000110010010" => q <= "00111010010100111010";
when "000110010011" => q <= "00111010110100110110";
when "000110010100" => q <= "00111011010100110010";
when "000110010101" => q <= "00111011100100101110";
when "000110010110" => q <= "00111100010100101010";
when "000110010111" => q <= "00111100110100100110";
when "000110011000" => q <= "00111101010100100001";
when "000110011001" => q <= "00111110000100011100";
when "000110011010" => q <= "00111110100100010111";
when "000110011011" => q <= "00111111010100010010";
when "000110011100" => q <= "01000000010100001011";
when "000110011101" => q <= "01000001000100000100";
when "000110011110" => q <= "01000010000011111100";
when "000110011111" => q <= "01000011000011110100";
when "000110100000" => q <= "01000100000011101010";
when "000110100001" => q <= "01000101000011100001";
when "000110100010" => q <= "01000101110011011000";
when "000110100011" => q <= "01000110100011010000";
when "000110100100" => q <= "01000110100011001011";
when "000110100101" => q <= "01000110000011001100";
when "000110100110" => q <= "01000100100011010101";
when "000110100111" => q <= "01000010000011101011";
when "000111000000" => q <= "00100111010011111011";
when "000111000001" => q <= "00101100110100110111";
when "000111000010" => q <= "00110000100101011100";
when "000111000011" => q <= "00110011010101110010";
when "000111000100" => q <= "00110101000101111011";
when "000111000101" => q <= "00110110000101111101";
when "000111000110" => q <= "00110110110101111010";
when "000111000111" => q <= "00110111000101110101";
when "000111001000" => q <= "00110111010101101110";
when "000111001001" => q <= "00110111010101100111";
when "000111001010" => q <= "00110111010101011111";
when "000111001011" => q <= "00110111010101011001";
when "000111001100" => q <= "00110111100101010011";
when "000111001101" => q <= "00110111100101001101";
when "000111001110" => q <= "00110111110101001001";
when "000111001111" => q <= "00111000000101000100";
when "000111010000" => q <= "00111000010101000000";
when "000111010001" => q <= "00111000110100111100";
when "000111010010" => q <= "00111001010100111000";
when "000111010011" => q <= "00111001100100110101";
when "000111010100" => q <= "00111010000100110001";
when "000111010101" => q <= "00111010100100101101";
when "000111010110" => q <= "00111011000100101001";
when "000111010111" => q <= "00111011100100100100";
when "000111011000" => q <= "00111100000100100000";
when "000111011001" => q <= "00111100100100011011";
when "000111011010" => q <= "00111101010100010110";
when "000111011011" => q <= "00111110000100010001";
when "000111011100" => q <= "00111110110100001011";
when "000111011101" => q <= "00111111100100000100";
when "000111011110" => q <= "01000000100011111100";
when "000111011111" => q <= "01000001010011110100";
when "000111100000" => q <= "01000010010011101011";
when "000111100001" => q <= "01000011010011100001";
when "000111100010" => q <= "01000100010011010111";
when "000111100011" => q <= "01000100110011001110";
when "000111100100" => q <= "01000101010011001000";
when "000111100101" => q <= "01000101000011000110";
when "000111100110" => q <= "01000100010011001011";
when "000111100111" => q <= "01000010010011011100";
when "001000000000" => q <= "00101001100100001111";
when "001000000001" => q <= "00101101110101000101";
when "001000000010" => q <= "00110000110101100101";
when "001000000011" => q <= "00110010110101110110";
when "001000000100" => q <= "00110100010101111101";
when "001000000101" => q <= "00110101000101111101";
when "001000000110" => q <= "00110101100101111001";
when "001000000111" => q <= "00110101110101110010";
when "001000001000" => q <= "00110101110101101011";
when "001000001001" => q <= "00110110000101100011";
when "001000001010" => q <= "00110110000101011100";
when "001000001011" => q <= "00110110000101010110";
when "001000001100" => q <= "00110110010101010000";
when "001000001101" => q <= "00110110010101001011";
when "001000001110" => q <= "00110110110101000110";
when "001000001111" => q <= "00110111000101000010";
when "001000010000" => q <= "00110111010100111110";
when "001000010001" => q <= "00110111110100111011";
when "001000010010" => q <= "00111000010100110111";
when "001000010011" => q <= "00111000100100110011";
when "001000010100" => q <= "00111001000100101111";
when "001000010101" => q <= "00111001100100101011";
when "001000010110" => q <= "00111010000100100111";
when "001000010111" => q <= "00111010100100100011";
when "001000011000" => q <= "00111011000100011111";
when "001000011001" => q <= "00111011100100011010";
when "001000011010" => q <= "00111100000100010101";
when "001000011011" => q <= "00111100110100010000";
when "001000011100" => q <= "00111101010100001010";
when "001000011101" => q <= "00111110000100000100";
when "001000011110" => q <= "00111110110011111100";
when "001000011111" => q <= "00111111110011110100";
when "001000100000" => q <= "01000000100011101011";
when "001000100001" => q <= "01000001100011100001";
when "001000100010" => q <= "01000010100011010111";
when "001000100011" => q <= "01000011010011001101";
when "001000100100" => q <= "01000011110011000101";
when "001000100101" => q <= "01000011110011000001";
when "001000100110" => q <= "01000011010011000100";
when "001000100111" => q <= "01000010010011010000";
when "001001000000" => q <= "00101010110100011110";
when "001001000001" => q <= "00101110010101001111";
when "001001000010" => q <= "00110000100101101011";
when "001001000011" => q <= "00110010000101111001";
when "001001000100" => q <= "00110011010101111110";
when "001001000101" => q <= "00110011110101111100";
when "001001000110" => q <= "00110100010101110111";
when "001001000111" => q <= "00110100100101110000";
when "001001001000" => q <= "00110100100101101000";
when "001001001001" => q <= "00110100100101100000";
when "001001001010" => q <= "00110100110101011001";
when "001001001011" => q <= "00110100110101010011";
when "001001001100" => q <= "00110101000101001101";
when "001001001101" => q <= "00110101010101001001";
when "001001001110" => q <= "00110101100101000100";
when "001001001111" => q <= "00110110000101000000";
when "001001010000" => q <= "00110110010100111101";
when "001001010001" => q <= "00110110110100111001";
when "001001010010" => q <= "00110111010100110101";
when "001001010011" => q <= "00110111110100110001";
when "001001010100" => q <= "00111000000100101110";
when "001001010101" => q <= "00111000100100101010";
when "001001010110" => q <= "00111001000100100110";
when "001001010111" => q <= "00111001100100100001";
when "001001011000" => q <= "00111010000100011101";
when "001001011001" => q <= "00111010100100011001";
when "001001011010" => q <= "00111011000100010100";
when "001001011011" => q <= "00111011100100001111";
when "001001011100" => q <= "00111100000100001001";
when "001001011101" => q <= "00111100110100000011";
when "001001011110" => q <= "00111101100011111100";
when "001001011111" => q <= "00111110010011110100";
when "001001100000" => q <= "00111111000011101011";
when "001001100001" => q <= "01000000000011100001";
when "001001100010" => q <= "01000000110011010110";
when "001001100011" => q <= "01000001100011001100";
when "001001100100" => q <= "01000010000011000011";
when "001001100101" => q <= "01000010010010111101";
when "001001100110" => q <= "01000010010010111110";
when "001001100111" => q <= "01000001100011000111";
when "001010000000" => q <= "00101011110100101010";
when "001010000001" => q <= "00101110010101010110";
when "001010000010" => q <= "00110000000101101111";
when "001010000011" => q <= "00110001010101111011";
when "001010000100" => q <= "00110010000101111110";
when "001010000101" => q <= "00110010100101111011";
when "001010000110" => q <= "00110011000101110101";
when "001010000111" => q <= "00110011000101101101";
when "001010001000" => q <= "00110011010101100101";
when "001010001001" => q <= "00110011100101011110";
when "001010001010" => q <= "00110011100101010111";
when "001010001011" => q <= "00110011110101010001";
when "001010001100" => q <= "00110100000101001011";
when "001010001101" => q <= "00110100010101000111";
when "001010001110" => q <= "00110100110101000010";
when "001010001111" => q <= "00110101000100111111";
when "001010010000" => q <= "00110101100100111011";
when "001010010001" => q <= "00110101110100110111";
when "001010010010" => q <= "00110110010100110100";
when "001010010011" => q <= "00110110110100110000";
when "001010010100" => q <= "00110111010100101100";
when "001010010101" => q <= "00110111100100101000";
when "001010010110" => q <= "00111000000100100100";
when "001010010111" => q <= "00111000100100100000";
when "001010011000" => q <= "00111001000100011100";
when "001010011001" => q <= "00111001010100010111";
when "001010011010" => q <= "00111001110100010011";
when "001010011011" => q <= "00111010010100001110";
when "001010011100" => q <= "00111010110100001000";
when "001010011101" => q <= "00111011100100000010";
when "001010011110" => q <= "00111100000011111011";
when "001010011111" => q <= "00111100110011110011";
when "001010100000" => q <= "00111101100011101010";
when "001010100001" => q <= "00111110010011100000";
when "001010100010" => q <= "00111111000011010110";
when "001010100011" => q <= "00111111110011001011";
when "001010100100" => q <= "01000000100011000001";
when "001010100101" => q <= "01000000110010111011";
when "001010100110" => q <= "01000000110010111001";
when "001010100111" => q <= "01000000100011000000";
when "001011000000" => q <= "00101100000100110010";
when "001011000001" => q <= "00101101110101011011";
when "001011000010" => q <= "00101111010101110010";
when "001011000011" => q <= "00110000010101111100";
when "001011000100" => q <= "00110000110101111101";
when "001011000101" => q <= "00110001010101111001";
when "001011000110" => q <= "00110001100101110011";
when "001011000111" => q <= "00110001110101101011";
when "001011001000" => q <= "00110010000101100011";
when "001011001001" => q <= "00110010010101011011";
when "001011001010" => q <= "00110010100101010100";
when "001011001011" => q <= "00110010110101001110";
when "001011001100" => q <= "00110011000101001001";
when "001011001101" => q <= "00110011010101000101";
when "001011001110" => q <= "00110011110101000001";
when "001011001111" => q <= "00110100000100111101";
when "001011010000" => q <= "00110100100100111001";
when "001011010001" => q <= "00110101000100110110";
when "001011010010" => q <= "00110101010100110010";
when "001011010011" => q <= "00110101110100101110";
when "001011010100" => q <= "00110110010100101011";
when "001011010101" => q <= "00110110110100100111";
when "001011010110" => q <= "00110111000100100010";
when "001011010111" => q <= "00110111100100011110";
when "001011011000" => q <= "00111000000100011010";
when "001011011001" => q <= "00111000010100010110";
when "001011011010" => q <= "00111000110100010001";
when "001011011011" => q <= "00111001010100001100";
when "001011011100" => q <= "00111001110100000111";
when "001011011101" => q <= "00111010010100000001";
when "001011011110" => q <= "00111010110011111010";
when "001011011111" => q <= "00111011100011110010";
when "001011100000" => q <= "00111100000011101010";
when "001011100001" => q <= "00111100110011100000";
when "001011100010" => q <= "00111101100011010101";
when "001011100011" => q <= "00111110010011001010";
when "001011100100" => q <= "00111110110011000000";
when "001011100101" => q <= "00111111010010111000";
when "001011100110" => q <= "00111111100010110101";
when "001011100111" => q <= "00111111010010111011";
when "001100000000" => q <= "00101100000100110111";
when "001100000001" => q <= "00101101010101011110";
when "001100000010" => q <= "00101110010101110011";
when "001100000011" => q <= "00101111000101111011";
when "001100000100" => q <= "00101111100101111100";
when "001100000101" => q <= "00110000000101111000";
when "001100000110" => q <= "00110000010101110001";
when "001100000111" => q <= "00110000110101101001";
when "001100001000" => q <= "00110001000101100001";
when "001100001001" => q <= "00110001010101011001";
when "001100001010" => q <= "00110001100101010010";
when "001100001011" => q <= "00110001110101001100";
when "001100001100" => q <= "00110010000101000111";
when "001100001101" => q <= "00110010100101000011";
when "001100001110" => q <= "00110010110100111111";
when "001100001111" => q <= "00110011010100111011";
when "001100010000" => q <= "00110011100100111000";
when "001100010001" => q <= "00110100000100110100";
when "001100010010" => q <= "00110100100100110001";
when "001100010011" => q <= "00110101000100101101";
when "001100010100" => q <= "00110101010100101001";
when "001100010101" => q <= "00110101110100100101";
when "001100010110" => q <= "00110110000100100001";
when "001100010111" => q <= "00110110100100011101";
when "001100011000" => q <= "00110111000100011000";
when "001100011001" => q <= "00110111010100010100";
when "001100011010" => q <= "00110111110100010000";
when "001100011011" => q <= "00111000010100001011";
when "001100011100" => q <= "00111000110100000110";
when "001100011101" => q <= "00111001000100000000";
when "001100011110" => q <= "00111001110011111001";
when "001100011111" => q <= "00111010010011110001";
when "001100100000" => q <= "00111010110011101001";
when "001100100001" => q <= "00111011010011011111";
when "001100100010" => q <= "00111100000011010100";
when "001100100011" => q <= "00111100100011001001";
when "001100100100" => q <= "00111101000010111110";
when "001100100101" => q <= "00111101100010110110";
when "001100100110" => q <= "00111101110010110011";
when "001100100111" => q <= "00111101110010110111";
when "001101000000" => q <= "00101100000100111001";
when "001101000001" => q <= "00101100110101011111";
when "001101000010" => q <= "00101101100101110011";
when "001101000011" => q <= "00101110000101111011";
when "001101000100" => q <= "00101110010101111011";
when "001101000101" => q <= "00101110110101110110";
when "001101000110" => q <= "00101111010101101111";
when "001101000111" => q <= "00101111100101100111";
when "001101001000" => q <= "00101111110101011111";
when "001101001001" => q <= "00110000010101010111";
when "001101001010" => q <= "00110000100101010000";
when "001101001011" => q <= "00110000110101001011";
when "001101001100" => q <= "00110001010101000110";
when "001101001101" => q <= "00110001100101000001";
when "001101001110" => q <= "00110010000100111110";
when "001101001111" => q <= "00110010010100111010";
when "001101010000" => q <= "00110010110100110110";
when "001101010001" => q <= "00110011000100110011";
when "001101010010" => q <= "00110011100100101111";
when "001101010011" => q <= "00110100000100101011";
when "001101010100" => q <= "00110100010100101000";
when "001101010101" => q <= "00110100110100100011";
when "001101010110" => q <= "00110101010100011111";
when "001101010111" => q <= "00110101100100011011";
when "001101011000" => q <= "00110110000100010111";
when "001101011001" => q <= "00110110010100010010";
when "001101011010" => q <= "00110110110100001110";
when "001101011011" => q <= "00110111010100001001";
when "001101011100" => q <= "00110111100100000100";
when "001101011101" => q <= "00111000000011111110";
when "001101011110" => q <= "00111000100011111000";
when "001101011111" => q <= "00111001000011110000";
when "001101100000" => q <= "00111001100011100111";
when "001101100001" => q <= "00111010000011011101";
when "001101100010" => q <= "00111010100011010011";
when "001101100011" => q <= "00111011000011000111";
when "001101100100" => q <= "00111011100010111101";
when "001101100101" => q <= "00111011110010110100";
when "001101100110" => q <= "00111100010010110000";
when "001101100111" => q <= "00111100100010110011";
when "001110000000" => q <= "00101011110100111010";
when "001110000001" => q <= "00101100000101011110";
when "001110000010" => q <= "00101100010101110010";
when "001110000011" => q <= "00101100110101111010";
when "001110000100" => q <= "00101101000101111010";
when "001110000101" => q <= "00101101100101110101";
when "001110000110" => q <= "00101110000101101110";
when "001110000111" => q <= "00101110010101100101";
when "001110001000" => q <= "00101110110101011101";
when "001110001001" => q <= "00101111000101010110";
when "001110001010" => q <= "00101111100101001111";
when "001110001011" => q <= "00101111110101001001";
when "001110001100" => q <= "00110000010101000100";
when "001110001101" => q <= "00110000110101000000";
when "001110001110" => q <= "00110001000100111100";
when "001110001111" => q <= "00110001100100111000";
when "001110010000" => q <= "00110001110100110101";
when "001110010001" => q <= "00110010010100110001";
when "001110010010" => q <= "00110010100100101110";
when "001110010011" => q <= "00110011000100101010";
when "001110010100" => q <= "00110011010100100110";
when "001110010101" => q <= "00110011110100100010";
when "001110010110" => q <= "00110100010100011110";
when "001110010111" => q <= "00110100100100011001";
when "001110011000" => q <= "00110101000100010101";
when "001110011001" => q <= "00110101010100010001";
when "001110011010" => q <= "00110101110100001100";
when "001110011011" => q <= "00110110000100001000";
when "001110011100" => q <= "00110110100100000010";
when "001110011101" => q <= "00110110110011111101";
when "001110011110" => q <= "00110111010011110110";
when "001110011111" => q <= "00110111110011101111";
when "001110100000" => q <= "00111000000011100110";
when "001110100001" => q <= "00111000100011011100";
when "001110100010" => q <= "00111001000011010001";
when "001110100011" => q <= "00111001010011000110";
when "001110100100" => q <= "00111001110010111011";
when "001110100101" => q <= "00111010010010110010";
when "001110100110" => q <= "00111010100010101110";
when "001110100111" => q <= "00111011000010110001";
when "001111000000" => q <= "00101011100100110111";
when "001111000001" => q <= "00101011010101011101";
when "001111000010" => q <= "00101011010101110000";
when "001111000011" => q <= "00101011100101111000";
when "001111000100" => q <= "00101011110101111000";
when "001111000101" => q <= "00101100010101110100";
when "001111000110" => q <= "00101100110101101100";
when "001111000111" => q <= "00101101000101100100";
when "001111001000" => q <= "00101101100101011100";
when "001111001001" => q <= "00101110000101010100";
when "001111001010" => q <= "00101110100101001110";
when "001111001011" => q <= "00101111000101001000";
when "001111001100" => q <= "00101111010101000011";
when "001111001101" => q <= "00101111110100111111";
when "001111001110" => q <= "00110000000100111011";
when "001111001111" => q <= "00110000100100110111";
when "001111010000" => q <= "00110001000100110100";
when "001111010001" => q <= "00110001010100110000";
when "001111010010" => q <= "00110001100100101100";
when "001111010011" => q <= "00110010000100101000";
when "001111010100" => q <= "00110010010100100100";
when "001111010101" => q <= "00110010110100100000";
when "001111010110" => q <= "00110011000100011100";
when "001111010111" => q <= "00110011100100011000";
when "001111011000" => q <= "00110100000100010100";
when "001111011001" => q <= "00110100010100001111";
when "001111011010" => q <= "00110100110100001011";
when "001111011011" => q <= "00110101000100000110";
when "001111011100" => q <= "00110101100100000001";
when "001111011101" => q <= "00110101110011111011";
when "001111011110" => q <= "00110110000011110100";
when "001111011111" => q <= "00110110100011101101";
when "001111100000" => q <= "00110110110011100100";
when "001111100001" => q <= "00110111000011011010";
when "001111100010" => q <= "00110111100011001111";
when "001111100011" => q <= "00110111110011000100";
when "001111100100" => q <= "00111000000010111001";
when "001111100101" => q <= "00111000100010110001";
when "001111100110" => q <= "00111001000010101100";
when "001111100111" => q <= "00111001010010110000";
when "010000000000" => q <= "00101011010100110011";
when "010000000001" => q <= "00101010110101011001";
when "010000000010" => q <= "00101010010101101110";
when "010000000011" => q <= "00101010010101110110";
when "010000000100" => q <= "00101010100101110111";
when "010000000101" => q <= "00101011000101110010";
when "010000000110" => q <= "00101011100101101011";
when "010000000111" => q <= "00101100000101100011";
when "010000001000" => q <= "00101100100101011011";
when "010000001001" => q <= "00101101000101010011";
when "010000001010" => q <= "00101101100101001101";
when "010000001011" => q <= "00101110000101000111";
when "010000001100" => q <= "00101110100101000010";
when "010000001101" => q <= "00101110110100111101";
when "010000001110" => q <= "00101111010100111001";
when "010000001111" => q <= "00101111100100110110";
when "010000010000" => q <= "00110000000100110010";
when "010000010001" => q <= "00110000010100101110";
when "010000010010" => q <= "00110000110100101011";
when "010000010011" => q <= "00110001000100100111";
when "010000010100" => q <= "00110001010100100011";
when "010000010101" => q <= "00110001110100011111";
when "010000010110" => q <= "00110010000100011011";
when "010000010111" => q <= "00110010100100010110";
when "010000011000" => q <= "00110010110100010010";
when "010000011001" => q <= "00110011010100001110";
when "010000011010" => q <= "00110011100100001001";
when "010000011011" => q <= "00110100000100000100";
when "010000011100" => q <= "00110100010011111111";
when "010000011101" => q <= "00110100100011111001";
when "010000011110" => q <= "00110101000011110010";
when "010000011111" => q <= "00110101010011101011";
when "010000100000" => q <= "00110101100011100010";
when "010000100001" => q <= "00110101110011011000";
when "010000100010" => q <= "00110110000011001101";
when "010000100011" => q <= "00110110000011000010";
when "010000100100" => q <= "00110110100010110111";
when "010000100101" => q <= "00110110110010101111";
when "010000100110" => q <= "00110111010010101011";
when "010000100111" => q <= "00111000000010101111";
when "010001000000" => q <= "00101011010100101011";
when "010001000001" => q <= "00101010000101010100";
when "010001000010" => q <= "00101001100101101010";
when "010001000011" => q <= "00101001010101110100";
when "010001000100" => q <= "00101001010101110101";
when "010001000101" => q <= "00101001110101110001";
when "010001000110" => q <= "00101010010101101011";
when "010001000111" => q <= "00101010110101100011";
when "010001001000" => q <= "00101011010101011010";
when "010001001001" => q <= "00101011110101010011";
when "010001001010" => q <= "00101100100101001100";
when "010001001011" => q <= "00101101000101000110";
when "010001001100" => q <= "00101101100101000001";
when "010001001101" => q <= "00101101110100111100";
when "010001001110" => q <= "00101110010100111000";
when "010001001111" => q <= "00101110110100110100";
when "010001010000" => q <= "00101111000100110001";
when "010001010001" => q <= "00101111010100101101";
when "010001010010" => q <= "00101111110100101001";
when "010001010011" => q <= "00110000000100100101";
when "010001010100" => q <= "00110000100100100001";
when "010001010101" => q <= "00110000110100011101";
when "010001010110" => q <= "00110001000100011001";
when "010001010111" => q <= "00110001100100010101";
when "010001011000" => q <= "00110001110100010000";
when "010001011001" => q <= "00110010010100001100";
when "010001011010" => q <= "00110010100100000111";
when "010001011011" => q <= "00110010110100000010";
when "010001011100" => q <= "00110011010011111101";
when "010001011101" => q <= "00110011100011110111";
when "010001011110" => q <= "00110011110011110000";
when "010001011111" => q <= "00110011110011101000";
when "010001100000" => q <= "00110100000011011111";
when "010001100001" => q <= "00110100010011010101";
when "010001100010" => q <= "00110100010011001010";
when "010001100011" => q <= "00110100100010111111";
when "010001100100" => q <= "00110100110010110101";
when "010001100101" => q <= "00110101000010101101";
when "010001100110" => q <= "00110101100010101010";
when "010001100111" => q <= "00110110100010110000";
when "010010000000" => q <= "00101011110100100001";
when "010010000001" => q <= "00101001110101001101";
when "010010000010" => q <= "00101000110101100101";
when "010010000011" => q <= "00101000010101110001";
when "010010000100" => q <= "00101000000101110011";
when "010010000101" => q <= "00101000010101110000";
when "010010000110" => q <= "00101000110101101010";
when "010010000111" => q <= "00101001100101100010";
when "010010001000" => q <= "00101010000101011010";
when "010010001001" => q <= "00101010110101010010";
when "010010001010" => q <= "00101011010101001011";
when "010010001011" => q <= "00101011110101000101";
when "010010001100" => q <= "00101100100101000000";
when "010010001101" => q <= "00101101000100111011";
when "010010001110" => q <= "00101101010100110111";
when "010010001111" => q <= "00101101110100110011";
when "010010010000" => q <= "00101110000100101111";
when "010010010001" => q <= "00101110100100101011";
when "010010010010" => q <= "00101110110100101000";
when "010010010011" => q <= "00101111000100100100";
when "010010010100" => q <= "00101111100100100000";
when "010010010101" => q <= "00101111110100011100";
when "010010010110" => q <= "00110000000100010111";
when "010010010111" => q <= "00110000100100010011";
when "010010011000" => q <= "00110000110100001111";
when "010010011001" => q <= "00110001000100001010";
when "010010011010" => q <= "00110001100100000110";
when "010010011011" => q <= "00110001110100000001";
when "010010011100" => q <= "00110010000011111011";
when "010010011101" => q <= "00110010010011110101";
when "010010011110" => q <= "00110010010011101110";
when "010010011111" => q <= "00110010100011100110";
when "010010100000" => q <= "00110010100011011101";
when "010010100001" => q <= "00110010100011010011";
when "010010100010" => q <= "00110010110011001000";
when "010010100011" => q <= "00110010110010111101";
when "010010100100" => q <= "00110011000010110011";
when "010010100101" => q <= "00110011100010101100";
when "010010100110" => q <= "00110100000010101010";
when "010010100111" => q <= "00110101000010110001";
when "010011000000" => q <= "00101100100100010100";
when "010011000001" => q <= "00101001110101000011";
when "010011000010" => q <= "00101000000101011111";
when "010011000011" => q <= "00100111010101101101";
when "010011000100" => q <= "00100111000101110001";
when "010011000101" => q <= "00100111000101101111";
when "010011000110" => q <= "00100111100101101001";
when "010011000111" => q <= "00101000000101100010";
when "010011001000" => q <= "00101000110101011010";
when "010011001001" => q <= "00101001100101010010";
when "010011001010" => q <= "00101010000101001011";
when "010011001011" => q <= "00101010110101000101";
when "010011001100" => q <= "00101011010100111111";
when "010011001101" => q <= "00101011110100111010";
when "010011001110" => q <= "00101100010100110110";
when "010011001111" => q <= "00101100110100110010";
when "010011010000" => q <= "00101101000100101110";
when "010011010001" => q <= "00101101100100101010";
when "010011010010" => q <= "00101101110100100110";
when "010011010011" => q <= "00101110000100100010";
when "010011010100" => q <= "00101110100100011110";
when "010011010101" => q <= "00101110110100011010";
when "010011010110" => q <= "00101111000100010110";
when "010011010111" => q <= "00101111100100010010";
when "010011011000" => q <= "00101111110100001101";
when "010011011001" => q <= "00110000000100001001";
when "010011011010" => q <= "00110000010100000100";
when "010011011011" => q <= "00110000100011111111";
when "010011011100" => q <= "00110000110011111001";
when "010011011101" => q <= "00110001000011110010";
when "010011011110" => q <= "00110001000011101011";
when "010011011111" => q <= "00110001000011100011";
when "010011100000" => q <= "00110001000011011010";
when "010011100001" => q <= "00110001000011001111";
when "010011100010" => q <= "00110001000011000101";
when "010011100011" => q <= "00110001000010111010";
when "010011100100" => q <= "00110001010010110001";
when "010011100101" => q <= "00110001110010101011";
when "010011100110" => q <= "00110010100010101011";
when "010011100111" => q <= "00110100000010110100";
when "010100000000" => q <= "00101101110100000010";
when "010100000001" => q <= "00101010000100110111";
when "010100000010" => q <= "00100111110101010111";
when "010100000011" => q <= "00100110100101100111";
when "010100000100" => q <= "00100101110101101110";
when "010100000101" => q <= "00100101110101101101";
when "010100000110" => q <= "00100110000101101001";
when "010100000111" => q <= "00100110100101100010";
when "010100001000" => q <= "00100111010101011010";
when "010100001001" => q <= "00101000000101010010";
when "010100001010" => q <= "00101000110101001011";
when "010100001011" => q <= "00101001100101000101";
when "010100001100" => q <= "00101010000100111111";
when "010100001101" => q <= "00101010110100111001";
when "010100001110" => q <= "00101011010100110101";
when "010100001111" => q <= "00101011110100110001";
when "010100010000" => q <= "00101100000100101100";
when "010100010001" => q <= "00101100100100101001";
when "010100010010" => q <= "00101100110100100101";
when "010100010011" => q <= "00101101000100100001";
when "010100010100" => q <= "00101101100100011101";
when "010100010101" => q <= "00101101110100011001";
when "010100010110" => q <= "00101110000100010100";
when "010100010111" => q <= "00101110010100010000";
when "010100011000" => q <= "00101110110100001100";
when "010100011001" => q <= "00101111000100000111";
when "010100011010" => q <= "00101111010100000010";
when "010100011011" => q <= "00101111010011111100";
when "010100011100" => q <= "00101111100011110110";
when "010100011101" => q <= "00101111100011110000";
when "010100011110" => q <= "00101111100011101000";
when "010100011111" => q <= "00101111100011100000";
when "010100100000" => q <= "00101111100011010110";
when "010100100001" => q <= "00101111010011001100";
when "010100100010" => q <= "00101111010011000010";
when "010100100011" => q <= "00101111010010111000";
when "010100100100" => q <= "00101111100010101111";
when "010100100101" => q <= "00110000010010101011";
when "010100100110" => q <= "00110001010010101101";
when "010100100111" => q <= "00110011010010111010";
when "010101000000" => q <= "00101111110011101100";
when "010101000001" => q <= "00101011000100100111";
when "010101000010" => q <= "00100111110101001100";
when "010101000011" => q <= "00100110000101100000";
when "010101000100" => q <= "00100101000101101001";
when "010101000101" => q <= "00100100100101101011";
when "010101000110" => q <= "00100100110101101000";
when "010101000111" => q <= "00100101010101100010";
when "010101001000" => q <= "00100101110101011010";
when "010101001001" => q <= "00100110100101010011";
when "010101001010" => q <= "00100111010101001011";
when "010101001011" => q <= "00101000000101000101";
when "010101001100" => q <= "00101000110100111111";
when "010101001101" => q <= "00101001100100111001";
when "010101001110" => q <= "00101010000100110100";
when "010101001111" => q <= "00101010100100110000";
when "010101010000" => q <= "00101011000100101011";
when "010101010001" => q <= "00101011010100100111";
when "010101010010" => q <= "00101011110100100011";
when "010101010011" => q <= "00101100000100011111";
when "010101010100" => q <= "00101100010100011011";
when "010101010101" => q <= "00101100110100010111";
when "010101010110" => q <= "00101101000100010011";
when "010101010111" => q <= "00101101010100001110";
when "010101011000" => q <= "00101101100100001010";
when "010101011001" => q <= "00101101110100000101";
when "010101011010" => q <= "00101101110100000000";
when "010101011011" => q <= "00101110000011111010";
when "010101011100" => q <= "00101110000011110100";
when "010101011101" => q <= "00101110000011101101";
when "010101011110" => q <= "00101110000011100101";
when "010101011111" => q <= "00101101110011011100";
when "010101100000" => q <= "00101101110011010011";
when "010101100001" => q <= "00101101100011001001";
when "010101100010" => q <= "00101101100010111111";
when "010101100011" => q <= "00101101100010110101";
when "010101100100" => q <= "00101110000010101110";
when "010101100101" => q <= "00101110110010101100";
when "010101100110" => q <= "00110000010010110001";
when "010101100111" => q <= "00110010110011000001";
when "010110000000" => q <= "00110011000011010000";
when "010110000001" => q <= "00101100110100010011";
when "010110000010" => q <= "00101000100100111110";
when "010110000011" => q <= "00100101110101010111";
when "010110000100" => q <= "00100100010101100011";
when "010110000101" => q <= "00100011100101100111";
when "010110000110" => q <= "00100011100101100110";
when "010110000111" => q <= "00100011110101100001";
when "010110001000" => q <= "00100100010101011011";
when "010110001001" => q <= "00100101000101010011";
when "010110001010" => q <= "00100101110101001100";
when "010110001011" => q <= "00100110100101000101";
when "010110001100" => q <= "00100111010100111111";
when "010110001101" => q <= "00101000000100111001";
when "010110001110" => q <= "00101000110100110100";
when "010110001111" => q <= "00101001010100101111";
when "010110010000" => q <= "00101001110100101010";
when "010110010001" => q <= "00101010000100100110";
when "010110010010" => q <= "00101010100100100010";
when "010110010011" => q <= "00101010110100011110";
when "010110010100" => q <= "00101011010100011010";
when "010110010101" => q <= "00101011100100010101";
when "010110010110" => q <= "00101011110100010001";
when "010110010111" => q <= "00101100000100001101";
when "010110011000" => q <= "00101100010100001000";
when "010110011001" => q <= "00101100010100000011";
when "010110011010" => q <= "00101100100011111101";
when "010110011011" => q <= "00101100100011110111";
when "010110011100" => q <= "00101100100011110001";
when "010110011101" => q <= "00101100010011101010";
when "010110011110" => q <= "00101100010011100001";
when "010110011111" => q <= "00101100000011011001";
when "010110100000" => q <= "00101011110011001111";
when "010110100001" => q <= "00101011100011000101";
when "010110100010" => q <= "00101011100010111100";
when "010110100011" => q <= "00101011110010110011";
when "010110100100" => q <= "00101100100010101110";
when "010110100101" => q <= "00101101110010101110";
when "010110100110" => q <= "00101111110010110111";
when "010110100111" => q <= "00110010110011001100";
when "010111000000" => q <= "00110111100010101110";
when "010111000001" => q <= "00101111110011111010";
when "010111000010" => q <= "00101010000100101100";
when "010111000011" => q <= "00100110010101001011";
when "010111000100" => q <= "00100100000101011011";
when "010111000101" => q <= "00100010110101100011";
when "010111000110" => q <= "00100010010101100011";
when "010111000111" => q <= "00100010010101100000";
when "010111001000" => q <= "00100010110101011010";
when "010111001001" => q <= "00100011010101010100";
when "010111001010" => q <= "00100100000101001101";
when "010111001011" => q <= "00100101000101000110";
when "010111001100" => q <= "00100101110100111111";
when "010111001101" => q <= "00100110100100111001";
when "010111001110" => q <= "00100111000100110100";
when "010111001111" => q <= "00100111110100101111";
when "010111010000" => q <= "00101000010100101010";
when "010111010001" => q <= "00101000110100100101";
when "010111010010" => q <= "00101001010100100001";
when "010111010011" => q <= "00101001100100011101";
when "010111010100" => q <= "00101001110100011000";
when "010111010101" => q <= "00101010000100010100";
when "010111010110" => q <= "00101010010100001111";
when "010111010111" => q <= "00101010100100001011";
when "010111011000" => q <= "00101010110100000110";
when "010111011001" => q <= "00101010110100000000";
when "010111011010" => q <= "00101010110011111011";
when "010111011011" => q <= "00101010110011110100";
when "010111011100" => q <= "00101010110011101110";
when "010111011101" => q <= "00101010100011100110";
when "010111011110" => q <= "00101010010011011110";
when "010111011111" => q <= "00101010000011010101";
when "010111100000" => q <= "00101001110011001011";
when "010111100001" => q <= "00101001110011000010";
when "010111100010" => q <= "00101001110010111001";
when "010111100011" => q <= "00101010010010110011";
when "010111100100" => q <= "00101011010010110000";
when "010111100101" => q <= "00101101000010110011";
when "010111100110" => q <= "00101111110011000000";
when "010111100111" => q <= "00110011110011011100";
when "011000000000" => q <= "00111110000010000011";
when "011000000001" => q <= "00110100000011011010";
when "011000000010" => q <= "00101100110100010101";
when "011000000011" => q <= "00100111110100111010";
when "011000000100" => q <= "00100100100101010001";
when "011000000101" => q <= "00100010100101011100";
when "011000000110" => q <= "00100001010101011111";
when "011000000111" => q <= "00100001000101011110";
when "011000001000" => q <= "00100001010101011010";
when "011000001001" => q <= "00100001110101010100";
when "011000001010" => q <= "00100010010101001101";
when "011000001011" => q <= "00100011000101000110";
when "011000001100" => q <= "00100100000101000000";
when "011000001101" => q <= "00100100110100111010";
when "011000001110" => q <= "00100101100100110100";
when "011000001111" => q <= "00100110000100101110";
when "011000010000" => q <= "00100110100100101001";
when "011000010001" => q <= "00100111000100100101";
when "011000010010" => q <= "00100111100100100000";
when "011000010011" => q <= "00101000000100011011";
when "011000010100" => q <= "00101000010100010111";
when "011000010101" => q <= "00101000100100010010";
when "011000010110" => q <= "00101000110100001101";
when "011000010111" => q <= "00101001000100001001";
when "011000011000" => q <= "00101001000100000011";
when "011000011001" => q <= "00101001000011111110";
when "011000011010" => q <= "00101001000011111000";
when "011000011011" => q <= "00101001000011110001";
when "011000011100" => q <= "00101000110011101010";
when "011000011101" => q <= "00101000100011100010";
when "011000011110" => q <= "00101000010011011010";
when "011000011111" => q <= "00101000000011010001";
when "011000100000" => q <= "00100111110011001000";
when "011000100001" => q <= "00100111110010111111";
when "011000100010" => q <= "00101000010010111000";
when "011000100011" => q <= "00101001000010110011";
when "011000100100" => q <= "00101010100010110011";
when "011000100101" => q <= "00101100110010111011";
when "011000100110" => q <= "00110000100011001101";
when "011000100111" => q <= "00110110000011110000";
when "011001000000" => q <= "01000110110001001101";
when "011001000001" => q <= "00111010010010110010";
when "011001000010" => q <= "00110001000011110111";
when "011001000011" => q <= "00101010010100100101";
when "011001000100" => q <= "00100101110101000010";
when "011001000101" => q <= "00100010110101010010";
when "011001000110" => q <= "00100001000101011001";
when "011001000111" => q <= "00100000000101011011";
when "011001001000" => q <= "00011111110101011000";
when "011001001001" => q <= "00100000000101010011";
when "011001001010" => q <= "00100000100101001101";
when "011001001011" => q <= "00100001010101000111";
when "011001001100" => q <= "00100010000101000000";
when "011001001101" => q <= "00100010110100111010";
when "011001001110" => q <= "00100011100100110100";
when "011001001111" => q <= "00100100000100101110";
when "011001010000" => q <= "00100100110100101001";
when "011001010001" => q <= "00100101010100100100";
when "011001010010" => q <= "00100101110100011111";
when "011001010011" => q <= "00100110010100011010";
when "011001010100" => q <= "00100110100100010101";
when "011001010101" => q <= "00100110110100010001";
when "011001010110" => q <= "00100111000100001100";
when "011001010111" => q <= "00100111000100000110";
when "011001011000" => q <= "00100111000100000001";
when "011001011001" => q <= "00100111000011111011";
when "011001011010" => q <= "00100111000011110101";
when "011001011011" => q <= "00100110110011101110";
when "011001011100" => q <= "00100110100011100110";
when "011001011101" => q <= "00100110010011011111";
when "011001011110" => q <= "00100110000011010110";
when "011001011111" => q <= "00100110000011001101";
when "011001100000" => q <= "00100110000011000101";
when "011001100001" => q <= "00100110000010111101";
when "011001100010" => q <= "00100110110010111000";
when "011001100011" => q <= "00101000000010110110";
when "011001100100" => q <= "00101010010010111010";
when "011001100101" => q <= "00101101110011000110";
when "011001100110" => q <= "00110010110011100000";
when "011001100111" => q <= "00111001110100001100";
when "011010000000" => q <= "01010010110000001100";
when "011010000001" => q <= "01000011000001111111";
when "011010000010" => q <= "00110111010011010001";
when "011010000011" => q <= "00101110100100001001";
when "011010000100" => q <= "00101000100100101110";
when "011010000101" => q <= "00100100000101000100";
when "011010000110" => q <= "00100001010101010000";
when "011010000111" => q <= "00011111110101010101";
when "011010001000" => q <= "00011111000101010101";
when "011010001001" => q <= "00011110110101010010";
when "011010001010" => q <= "00011111000101001101";
when "011010001011" => q <= "00011111010101000111";
when "011010001100" => q <= "00100000000101000001";
when "011010001101" => q <= "00100000110100111010";
when "011010001110" => q <= "00100001010100110100";
when "011010001111" => q <= "00100010000100101110";
when "011010010000" => q <= "00100010110100101001";
when "011010010001" => q <= "00100011010100100011";
when "011010010010" => q <= "00100011110100011110";
when "011010010011" => q <= "00100100000100011001";
when "011010010100" => q <= "00100100100100010100";
when "011010010101" => q <= "00100100110100001111";
when "011010010110" => q <= "00100100110100001010";
when "011010010111" => q <= "00100101000100000100";
when "011010011000" => q <= "00100101000011111110";
when "011010011001" => q <= "00100100110011111000";
when "011010011010" => q <= "00100100110011110001";
when "011010011011" => q <= "00100100100011101010";
when "011010011100" => q <= "00100100010011100011";
when "011010011101" => q <= "00100100000011011011";
when "011010011110" => q <= "00100100000011010011";
when "011010011111" => q <= "00100100000011001011";
when "011010100000" => q <= "00100100010011000011";
when "011010100001" => q <= "00100100110010111101";
when "011010100010" => q <= "00100110000010111010";
when "011010100011" => q <= "00101000000010111100";
when "011010100100" => q <= "00101011000011000100";
when "011010100101" => q <= "00101111110011010111";
when "011010100110" => q <= "00110110100011111001";
when "011010100111" => q <= "00111111100100110000";
when "011011000000" => q <= "01100010100000000000";
when "011011000001" => q <= "01001111010001000001";
when "011011000010" => q <= "01000000010010100010";
when "011011000011" => q <= "00110101000011100110";
when "011011000100" => q <= "00101100110100010100";
when "011011000101" => q <= "00100111000100110010";
when "011011000110" => q <= "00100010110101000011";
when "011011000111" => q <= "00100000010101001100";
when "011011001000" => q <= "00011110100101010000";
when "011011001001" => q <= "00011101110101001111";
when "011011001010" => q <= "00011101100101001011";
when "011011001011" => q <= "00011101110101000110";
when "011011001100" => q <= "00011110000101000001";
when "011011001101" => q <= "00011110100100111011";
when "011011001110" => q <= "00011111010100110101";
when "011011001111" => q <= "00011111110100101111";
when "011011010000" => q <= "00100000010100101001";
when "011011010001" => q <= "00100001000100100011";
when "011011010010" => q <= "00100001010100011101";
when "011011010011" => q <= "00100001110100011000";
when "011011010100" => q <= "00100010000100010011";
when "011011010101" => q <= "00100010010100001101";
when "011011010110" => q <= "00100010100100000111";
when "011011010111" => q <= "00100010100100000010";
when "011011011000" => q <= "00100010100011111100";
when "011011011001" => q <= "00100010100011110101";
when "011011011010" => q <= "00100010010011101110";
when "011011011011" => q <= "00100010010011100111";
when "011011011100" => q <= "00100010000011011111";
when "011011011101" => q <= "00100010000011011000";
when "011011011110" => q <= "00100010000011010000";
when "011011011111" => q <= "00100010010011001001";
when "011011100000" => q <= "00100010110011000011";
when "011011100001" => q <= "00100100000010111111";
when "011011100010" => q <= "00100110000010111111";
when "011011100011" => q <= "00101001000011000101";
when "011011100100" => q <= "00101101100011010100";
when "011011100101" => q <= "00110011110011101111";
when "011011100110" => q <= "00111100100100011011";
when "011011100111" => q <= "01001000010101011110";
when "011100000000" => q <= "01110000000000000000";
when "011100000001" => q <= "01011111100000000000";
when "011100000010" => q <= "01001101000001100110";
when "011100000011" => q <= "00111110110010111000";
when "011100000100" => q <= "00110011110011110010";
when "011100000101" => q <= "00101011110100011000";
when "011100000110" => q <= "00100110000100110001";
when "011100000111" => q <= "00100010000101000000";
when "011100001000" => q <= "00011111010101000111";
when "011100001001" => q <= "00011101110101001001";
when "011100001010" => q <= "00011100110101001000";
when "011100001011" => q <= "00011100100101000100";
when "011100001100" => q <= "00011100100101000000";
when "011100001101" => q <= "00011100110100111010";
when "011100001110" => q <= "00011101000100110100";
when "011100001111" => q <= "00011101100100101110";
when "011100010000" => q <= "00011110000100101000";
when "011100010001" => q <= "00011110100100100011";
when "011100010010" => q <= "00011111000100011101";
when "011100010011" => q <= "00011111010100010111";
when "011100010100" => q <= "00011111100100010001";
when "011100010101" => q <= "00011111110100001011";
when "011100010110" => q <= "00100000000100000101";
when "011100010111" => q <= "00100000000011111111";
when "011100011000" => q <= "00100000000011111001";
when "011100011001" => q <= "00100000000011110010";
when "011100011010" => q <= "00100000000011101011";
when "011100011011" => q <= "00100000000011100100";
when "011100011100" => q <= "00100000000011011101";
when "011100011101" => q <= "00100000000011010101";
when "011100011110" => q <= "00100000100011001111";
when "011100011111" => q <= "00100001010011001001";
when "011100100000" => q <= "00100010100011000101";
when "011100100001" => q <= "00100100010011000101";
when "011100100010" => q <= "00100111100011001001";
when "011100100011" => q <= "00101011110011010101";
when "011100100100" => q <= "00110010000011101011";
when "011100100101" => q <= "00111010010100001111";
when "011100100110" => q <= "01000101110101001000";
when "011100100111" => q <= "01010100110110011010";
when "011101000000" => q <= "01110000000000000000";
when "011101000001" => q <= "01110000000000000000";
when "011101000010" => q <= "01011110010000011011";
when "011101000011" => q <= "01001100000001111110";
when "011101000100" => q <= "00111110000011000101";
when "011101000101" => q <= "00110011100011110111";
when "011101000110" => q <= "00101011100100011000";
when "011101000111" => q <= "00100101110100101110";
when "011101001000" => q <= "00100001110100111010";
when "011101001001" => q <= "00011110110101000000";
when "011101001010" => q <= "00011101000101000010";
when "011101001011" => q <= "00011100000101000000";
when "011101001100" => q <= "00011011100100111101";
when "011101001101" => q <= "00011011010100111001";
when "011101001110" => q <= "00011011010100110011";
when "011101001111" => q <= "00011011100100101110";
when "011101010000" => q <= "00011100000100101000";
when "011101010001" => q <= "00011100010100100010";
when "011101010010" => q <= "00011100100100011100";
when "011101010011" => q <= "00011100110100010110";
when "011101010100" => q <= "00011101010100010000";
when "011101010101" => q <= "00011101010100001010";
when "011101010110" => q <= "00011101100100000011";
when "011101010111" => q <= "00011101100011111101";
when "011101011000" => q <= "00011101110011110110";
when "011101011001" => q <= "00011101110011110000";
when "011101011010" => q <= "00011101110011101001";
when "011101011011" => q <= "00011110000011100010";
when "011101011100" => q <= "00011110010011011011";
when "011101011101" => q <= "00011110110011010101";
when "011101011110" => q <= "00011111110011001111";
when "011101011111" => q <= "00100001000011001100";
when "011101100000" => q <= "00100011010011001011";
when "011101100001" => q <= "00100110010011001110";
when "011101100010" => q <= "00101010110011011000";
when "011101100011" => q <= "00110000110011101011";
when "011101100100" => q <= "00111001010100001010";
when "011101100101" => q <= "01000100010100111011";
when "011101100110" => q <= "01010011000110000001";
when "011101100111" => q <= "01100110000111000000";

      when others => q <=   "00000000000000000000";
    end case;
  end process;

end rtl;

