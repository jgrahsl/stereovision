../sim_pkg.vhd