
library ieee;
use ieee.std_logic_1164.all;
library work;
use work.cam_pkg.all;

entity romdata is
  generic (ADR_BITS  : integer;
           DATA_BITS : integer);             -- for compatibility
  port (
    clk : in  std_logic;
    a   : in  std_logic_vector(ADR_BITS-1 downto 0);
    q   : out std_logic_vector(DATA_BITS-1 downto 0));
end romdata;

architecture rtl of romdata is
    ATTRIBUTE ram_extract: string;
    ATTRIBUTE ram_extract OF q: SIGNAL IS "yes";
    ATTRIBUTE ram_style: string;
    ATTRIBUTE ram_style OF q: SIGNAL IS "block";
  
  signal areg : std_logic_vector((GRIDX_BITS+GRIDY_BITS-1) downto 0);  -- GRIDX+GRIDY-1
begin

  process(clk)
  begin
    if rising_edge(clk) then
      areg <= a(areg'high downto areg'low);
    end if;
  end process;

  process(areg)
  begin
    case areg is
      -- GRIDY+GRIDX --    REFY+REFX

when "000000000000" => q <= "00000000000000000000";
when "000000000001" => q <= "00000000000000000000";
when "000000000010" => q <= "00000000000000000000";
when "000000000011" => q <= "00000000000000110101";
when "000000000100" => q <= "00000000000001110001";
when "000000000101" => q <= "00000101100010000000";
when "000000000110" => q <= "00001100000010000000";
when "000000000111" => q <= "00010000110010000000";
when "000000001000" => q <= "00010100100010000000";
when "000000001001" => q <= "00010111000010000000";
when "000000001010" => q <= "00011000110010000000";
when "000000001011" => q <= "00011001110010000000";
when "000000001100" => q <= "00011010110010000000";
when "000000001101" => q <= "00011011010010000000";
when "000000001110" => q <= "00011011110010000000";
when "000000001111" => q <= "00011100000010000000";
when "000000010000" => q <= "00011100010010000000";
when "000000010001" => q <= "00011100110010000000";
when "000000010010" => q <= "00011101000010000000";
when "000000010011" => q <= "00011101100010000000";
when "000000010100" => q <= "00011110000010000000";
when "000000010101" => q <= "00011110100010000000";
when "000000010110" => q <= "00011111010010000000";
when "000000010111" => q <= "00100000000010000000";
when "000000011000" => q <= "00100000000010000000";
when "000000011001" => q <= "00100000000010000000";
when "000000011010" => q <= "00100000000001111001";
when "000000011011" => q <= "00100000000001110010";
when "000000011100" => q <= "00100000000001101100";
when "000000011101" => q <= "00100000000001100101";
when "000000011110" => q <= "00100000000001011111";
when "000000011111" => q <= "00100000000001011010";
when "000000100000" => q <= "00100000000001010110";
when "000000100001" => q <= "00100000000001010111";
when "000000100010" => q <= "00100000000001011100";
when "000000100011" => q <= "00011100100001101000";
when "000000100100" => q <= "00010110110001111111";
when "000000100101" => q <= "00001110110010000000";
when "000000100110" => q <= "00000011100010000000";
when "000000100111" => q <= "00000000000010000000";
when "000001000000" => q <= "00000000000000000000";
when "000001000001" => q <= "00000000000000000000";
when "000001000010" => q <= "00000000000000011100";
when "000001000011" => q <= "00000000000001100010";
when "000001000100" => q <= "00000100000010000000";
when "000001000101" => q <= "00001010100010000000";
when "000001000110" => q <= "00001111100010000000";
when "000001000111" => q <= "00010011000010000000";
when "000001001000" => q <= "00010101100010000000";
when "000001001001" => q <= "00010111000010000000";
when "000001001010" => q <= "00011000010010000000";
when "000001001011" => q <= "00011000110010000000";
when "000001001100" => q <= "00011001010010000000";
when "000001001101" => q <= "00011001100010000000";
when "000001001110" => q <= "00011001110010000000";
when "000001001111" => q <= "00011010000010000000";
when "000001010000" => q <= "00011010010010000000";
when "000001010001" => q <= "00011010100010000000";
when "000001010010" => q <= "00011010110010000000";
when "000001010011" => q <= "00011011010010000000";
when "000001010100" => q <= "00011011110010000000";
when "000001010101" => q <= "00011100010010000000";
when "000001010110" => q <= "00011100110010000000";
when "000001010111" => q <= "00011101100010000000";
when "000001011000" => q <= "00011110010010000000";
when "000001011001" => q <= "00011111010001111111";
when "000001011010" => q <= "00100000000001111001";
when "000001011011" => q <= "00100000000001110010";
when "000001011100" => q <= "00100000000001101011";
when "000001011101" => q <= "00100000000001100100";
when "000001011110" => q <= "00100000000001011100";
when "000001011111" => q <= "00100000000001010110";
when "000001100000" => q <= "00100000000001010000";
when "000001100001" => q <= "00100000000001001101";
when "000001100010" => q <= "00100000000001001110";
when "000001100011" => q <= "00011111110001010101";
when "000001100100" => q <= "00011011110001100100";
when "000001100101" => q <= "00010110000010000000";
when "000001100110" => q <= "00001101100010000000";
when "000001100111" => q <= "00000001110010000000";
when "000010000000" => q <= "00000000000000000000";
when "000010000001" => q <= "00000000000000000000";
when "000010000010" => q <= "00000000000001001011";
when "000010000011" => q <= "00000001110010000000";
when "000010000100" => q <= "00001000100010000000";
when "000010000101" => q <= "00001101110010000000";
when "000010000110" => q <= "00010001010010000000";
when "000010000111" => q <= "00010011110010000000";
when "000010001000" => q <= "00010101010010000000";
when "000010001001" => q <= "00010110100010000000";
when "000010001010" => q <= "00010111000010000000";
when "000010001011" => q <= "00010111100010000000";
when "000010001100" => q <= "00010111100010000000";
when "000010001101" => q <= "00010111110010000000";
when "000010001110" => q <= "00010111110010000000";
when "000010001111" => q <= "00011000000010000000";
when "000010010000" => q <= "00011000010010000000";
when "000010010001" => q <= "00011000010010000000";
when "000010010010" => q <= "00011000110010000000";
when "000010010011" => q <= "00011001000010000000";
when "000010010100" => q <= "00011001100010000000";
when "000010010101" => q <= "00011010000010000000";
when "000010010110" => q <= "00011010110010000000";
when "000010010111" => q <= "00011011010010000000";
when "000010011000" => q <= "00011100010010000000";
when "000010011001" => q <= "00011101000001111111";
when "000010011010" => q <= "00011110000001111001";
when "000010011011" => q <= "00011110110001110010";
when "000010011100" => q <= "00011111110001101011";
when "000010011101" => q <= "00100000000001100011";
when "000010011110" => q <= "00100000000001011011";
when "000010011111" => q <= "00100000000001010100";
when "000010100000" => q <= "00100000000001001101";
when "000010100001" => q <= "00100000000001001000";
when "000010100010" => q <= "00100000000001000101";
when "000010100011" => q <= "00100000000001000111";
when "000010100100" => q <= "00011110110001010001";
when "000010100101" => q <= "00011010100001100100";
when "000010100110" => q <= "00010100010010000000";
when "000010100111" => q <= "00001011010010000000";
when "000011000000" => q <= "00000000000000000000";
when "000011000001" => q <= "00000000000000101000";
when "000011000010" => q <= "00000000000001101111";
when "000011000011" => q <= "00000110010010000000";
when "000011000100" => q <= "00001011100010000000";
when "000011000101" => q <= "00001111010010000000";
when "000011000110" => q <= "00010001110010000000";
when "000011000111" => q <= "00010011100010000000";
when "000011001000" => q <= "00010100110010000000";
when "000011001001" => q <= "00010101010010000000";
when "000011001010" => q <= "00010101100010000000";
when "000011001011" => q <= "00010101110010000000";
when "000011001100" => q <= "00010101110010000000";
when "000011001101" => q <= "00010101110010000000";
when "000011001110" => q <= "00010110000010000000";
when "000011001111" => q <= "00010110000010000000";
when "000011010000" => q <= "00010110010010000000";
when "000011010001" => q <= "00010110100010000000";
when "000011010010" => q <= "00010110110010000000";
when "000011010011" => q <= "00010111000010000000";
when "000011010100" => q <= "00010111100010000000";
when "000011010101" => q <= "00011000000010000000";
when "000011010110" => q <= "00011000110010000000";
when "000011010111" => q <= "00011001010010000000";
when "000011011000" => q <= "00011010000010000000";
when "000011011001" => q <= "00011011000001111110";
when "000011011010" => q <= "00011011110001111000";
when "000011011011" => q <= "00011100110001110010";
when "000011011100" => q <= "00011101110001101011";
when "000011011101" => q <= "00011110110001100011";
when "000011011110" => q <= "00011111110001011011";
when "000011011111" => q <= "00100000000001010011";
when "000011100000" => q <= "00100000000001001011";
when "000011100001" => q <= "00100000000001000100";
when "000011100010" => q <= "00100000000000111111";
when "000011100011" => q <= "00100000000000111110";
when "000011100100" => q <= "00100000000001000010";
when "000011100101" => q <= "00011101010001010000";
when "000011100110" => q <= "00011000100001101010";
when "000011100111" => q <= "00010001110010000000";
when "000100000000" => q <= "00000000000000000000";
when "000100000001" => q <= "00000000000001001110";
when "000100000010" => q <= "00000011010010000000";
when "000100000011" => q <= "00001001000010000000";
when "000100000100" => q <= "00001101000010000000";
when "000100000101" => q <= "00001111110010000000";
when "000100000110" => q <= "00010001110010000000";
when "000100000111" => q <= "00010010110010000000";
when "000100001000" => q <= "00010011100010000000";
when "000100001001" => q <= "00010011110010000000";
when "000100001010" => q <= "00010100000010000000";
when "000100001011" => q <= "00010100000010000000";
when "000100001100" => q <= "00010100000010000000";
when "000100001101" => q <= "00010100000010000000";
when "000100001110" => q <= "00010100000010000000";
when "000100001111" => q <= "00010100010010000000";
when "000100010000" => q <= "00010100100010000000";
when "000100010001" => q <= "00010100110010000000";
when "000100010010" => q <= "00010101000010000000";
when "000100010011" => q <= "00010101100010000000";
when "000100010100" => q <= "00010101110010000000";
when "000100010101" => q <= "00010110010010000000";
when "000100010110" => q <= "00010111000010000000";
when "000100010111" => q <= "00010111100010000000";
when "000100011000" => q <= "00011000010010000000";
when "000100011001" => q <= "00011001000001111110";
when "000100011010" => q <= "00011001110001111000";
when "000100011011" => q <= "00011010110001110010";
when "000100011100" => q <= "00011011110001101011";
when "000100011101" => q <= "00011100110001100100";
when "000100011110" => q <= "00011101110001011100";
when "000100011111" => q <= "00011110110001010011";
when "000100100000" => q <= "00011111110001001010";
when "000100100001" => q <= "00100000000001000010";
when "000100100010" => q <= "00100000000000111011";
when "000100100011" => q <= "00100000000000110111";
when "000100100100" => q <= "00100000000000111000";
when "000100100101" => q <= "00011110010001000000";
when "000100100110" => q <= "00011011000001010011";
when "000100100111" => q <= "00010110000001110110";
when "000101000000" => q <= "00000000000000011111";
when "000101000001" => q <= "00000000000001101101";
when "000101000010" => q <= "00000110000010000000";
when "000101000011" => q <= "00001010100010000000";
when "000101000100" => q <= "00001101100010000000";
when "000101000101" => q <= "00001111110010000000";
when "000101000110" => q <= "00010001000010000000";
when "000101000111" => q <= "00010001110010000000";
when "000101001000" => q <= "00010010000010000000";
when "000101001001" => q <= "00010010010010000000";
when "000101001010" => q <= "00010010010010000000";
when "000101001011" => q <= "00010010010010000000";
when "000101001100" => q <= "00010010010010000000";
when "000101001101" => q <= "00010010010010000000";
when "000101001110" => q <= "00010010100010000000";
when "000101001111" => q <= "00010010110010000000";
when "000101010000" => q <= "00010010110010000000";
when "000101010001" => q <= "00010011010010000000";
when "000101010010" => q <= "00010011100010000000";
when "000101010011" => q <= "00010100000010000000";
when "000101010100" => q <= "00010100100010000000";
when "000101010101" => q <= "00010101000010000000";
when "000101010110" => q <= "00010101100010000000";
when "000101010111" => q <= "00010110000010000000";
when "000101011000" => q <= "00010110110010000000";
when "000101011001" => q <= "00010111010001111101";
when "000101011010" => q <= "00011000000001111000";
when "000101011011" => q <= "00011001000001110010";
when "000101011100" => q <= "00011001110001101011";
when "000101011101" => q <= "00011010110001100100";
when "000101011110" => q <= "00011011110001011100";
when "000101011111" => q <= "00011101000001010011";
when "000101100000" => q <= "00011110000001001010";
when "000101100001" => q <= "00011110110001000001";
when "000101100010" => q <= "00011111100000111001";
when "000101100011" => q <= "00011111110000110011";
when "000101100100" => q <= "00011111100000110001";
when "000101100101" => q <= "00011110100000110101";
when "000101100110" => q <= "00011100010001000010";
when "000101100111" => q <= "00011000100001011110";
when "000110000000" => q <= "00000000000001000001";
when "000110000001" => q <= "00000010110010000000";
when "000110000010" => q <= "00000111110010000000";
when "000110000011" => q <= "00001011010010000000";
when "000110000100" => q <= "00001101100010000000";
when "000110000101" => q <= "00001111000010000000";
when "000110000110" => q <= "00010000000010000000";
when "000110000111" => q <= "00010000100010000000";
when "000110001000" => q <= "00010000110010000000";
when "000110001001" => q <= "00010000110010000000";
when "000110001010" => q <= "00010000110010000000";
when "000110001011" => q <= "00010000110010000000";
when "000110001100" => q <= "00010000110010000000";
when "000110001101" => q <= "00010001000010000000";
when "000110001110" => q <= "00010001000010000000";
when "000110001111" => q <= "00010001010010000000";
when "000110010000" => q <= "00010001100010000000";
when "000110010001" => q <= "00010001110010000000";
when "000110010010" => q <= "00010010010010000000";
when "000110010011" => q <= "00010010110010000000";
when "000110010100" => q <= "00010011010010000000";
when "000110010101" => q <= "00010011100010000000";
when "000110010110" => q <= "00010100010010000000";
when "000110010111" => q <= "00010100110010000000";
when "000110011000" => q <= "00010101010010000000";
when "000110011001" => q <= "00010110000001111100";
when "000110011010" => q <= "00010110100001110111";
when "000110011011" => q <= "00010111010001110010";
when "000110011100" => q <= "00011000010001101011";
when "000110011101" => q <= "00011001000001100100";
when "000110011110" => q <= "00011010000001011100";
when "000110011111" => q <= "00011011000001010100";
when "000110100000" => q <= "00011100000001001010";
when "000110100001" => q <= "00011101000001000001";
when "000110100010" => q <= "00011101110000111000";
when "000110100011" => q <= "00011110100000110000";
when "000110100100" => q <= "00011110100000101011";
when "000110100101" => q <= "00011110000000101100";
when "000110100110" => q <= "00011100100000110101";
when "000110100111" => q <= "00011010000001001011";
when "000111000000" => q <= "00000000000001011011";
when "000111000001" => q <= "00000100110010000000";
when "000111000010" => q <= "00001000100010000000";
when "000111000011" => q <= "00001011010010000000";
when "000111000100" => q <= "00001101000010000000";
when "000111000101" => q <= "00001110000010000000";
when "000111000110" => q <= "00001110110010000000";
when "000111000111" => q <= "00001111000010000000";
when "000111001000" => q <= "00001111010010000000";
when "000111001001" => q <= "00001111010010000000";
when "000111001010" => q <= "00001111010010000000";
when "000111001011" => q <= "00001111010010000000";
when "000111001100" => q <= "00001111100010000000";
when "000111001101" => q <= "00001111100010000000";
when "000111001110" => q <= "00001111110010000000";
when "000111001111" => q <= "00010000000010000000";
when "000111010000" => q <= "00010000010010000000";
when "000111010001" => q <= "00010000110010000000";
when "000111010010" => q <= "00010001010010000000";
when "000111010011" => q <= "00010001100010000000";
when "000111010100" => q <= "00010010000010000000";
when "000111010101" => q <= "00010010100010000000";
when "000111010110" => q <= "00010011000010000000";
when "000111010111" => q <= "00010011100010000000";
when "000111011000" => q <= "00010100000010000000";
when "000111011001" => q <= "00010100100001111011";
when "000111011010" => q <= "00010101010001110110";
when "000111011011" => q <= "00010110000001110001";
when "000111011100" => q <= "00010110110001101011";
when "000111011101" => q <= "00010111100001100100";
when "000111011110" => q <= "00011000100001011100";
when "000111011111" => q <= "00011001010001010100";
when "000111100000" => q <= "00011010010001001011";
when "000111100001" => q <= "00011011010001000001";
when "000111100010" => q <= "00011100010000110111";
when "000111100011" => q <= "00011100110000101110";
when "000111100100" => q <= "00011101010000101000";
when "000111100101" => q <= "00011101000000100110";
when "000111100110" => q <= "00011100010000101011";
when "000111100111" => q <= "00011010010000111100";
when "001000000000" => q <= "00000001100001101111";
when "001000000001" => q <= "00000101110010000000";
when "001000000010" => q <= "00001000110010000000";
when "001000000011" => q <= "00001010110010000000";
when "001000000100" => q <= "00001100010010000000";
when "001000000101" => q <= "00001101000010000000";
when "001000000110" => q <= "00001101100010000000";
when "001000000111" => q <= "00001101110010000000";
when "001000001000" => q <= "00001101110010000000";
when "001000001001" => q <= "00001110000010000000";
when "001000001010" => q <= "00001110000010000000";
when "001000001011" => q <= "00001110000010000000";
when "001000001100" => q <= "00001110010010000000";
when "001000001101" => q <= "00001110010010000000";
when "001000001110" => q <= "00001110110010000000";
when "001000001111" => q <= "00001111000010000000";
when "001000010000" => q <= "00001111010010000000";
when "001000010001" => q <= "00001111110010000000";
when "001000010010" => q <= "00010000010010000000";
when "001000010011" => q <= "00010000100010000000";
when "001000010100" => q <= "00010001000010000000";
when "001000010101" => q <= "00010001100010000000";
when "001000010110" => q <= "00010010000010000000";
when "001000010111" => q <= "00010010100010000000";
when "001000011000" => q <= "00010011000001111111";
when "001000011001" => q <= "00010011100001111010";
when "001000011010" => q <= "00010100000001110101";
when "001000011011" => q <= "00010100110001110000";
when "001000011100" => q <= "00010101010001101010";
when "001000011101" => q <= "00010110000001100100";
when "001000011110" => q <= "00010110110001011100";
when "001000011111" => q <= "00010111110001010100";
when "001000100000" => q <= "00011000100001001011";
when "001000100001" => q <= "00011001100001000001";
when "001000100010" => q <= "00011010100000110111";
when "001000100011" => q <= "00011011010000101101";
when "001000100100" => q <= "00011011110000100101";
when "001000100101" => q <= "00011011110000100001";
when "001000100110" => q <= "00011011010000100100";
when "001000100111" => q <= "00011010010000110000";
when "001001000000" => q <= "00000010110001111110";
when "001001000001" => q <= "00000110010010000000";
when "001001000010" => q <= "00001000100010000000";
when "001001000011" => q <= "00001010000010000000";
when "001001000100" => q <= "00001011010010000000";
when "001001000101" => q <= "00001011110010000000";
when "001001000110" => q <= "00001100010010000000";
when "001001000111" => q <= "00001100100010000000";
when "001001001000" => q <= "00001100100010000000";
when "001001001001" => q <= "00001100100010000000";
when "001001001010" => q <= "00001100110010000000";
when "001001001011" => q <= "00001100110010000000";
when "001001001100" => q <= "00001101000010000000";
when "001001001101" => q <= "00001101010010000000";
when "001001001110" => q <= "00001101100010000000";
when "001001001111" => q <= "00001110000010000000";
when "001001010000" => q <= "00001110010010000000";
when "001001010001" => q <= "00001110110010000000";
when "001001010010" => q <= "00001111010010000000";
when "001001010011" => q <= "00001111110010000000";
when "001001010100" => q <= "00010000000010000000";
when "001001010101" => q <= "00010000100010000000";
when "001001010110" => q <= "00010001000010000000";
when "001001010111" => q <= "00010001100010000000";
when "001001011000" => q <= "00010010000001111101";
when "001001011001" => q <= "00010010100001111001";
when "001001011010" => q <= "00010011000001110100";
when "001001011011" => q <= "00010011100001101111";
when "001001011100" => q <= "00010100000001101001";
when "001001011101" => q <= "00010100110001100011";
when "001001011110" => q <= "00010101100001011100";
when "001001011111" => q <= "00010110010001010100";
when "001001100000" => q <= "00010111000001001011";
when "001001100001" => q <= "00011000000001000001";
when "001001100010" => q <= "00011000110000110110";
when "001001100011" => q <= "00011001100000101100";
when "001001100100" => q <= "00011010000000100011";
when "001001100101" => q <= "00011010010000011101";
when "001001100110" => q <= "00011010010000011110";
when "001001100111" => q <= "00011001100000100111";
when "001010000000" => q <= "00000011110010000000";
when "001010000001" => q <= "00000110010010000000";
when "001010000010" => q <= "00001000000010000000";
when "001010000011" => q <= "00001001010010000000";
when "001010000100" => q <= "00001010000010000000";
when "001010000101" => q <= "00001010100010000000";
when "001010000110" => q <= "00001011000010000000";
when "001010000111" => q <= "00001011000010000000";
when "001010001000" => q <= "00001011010010000000";
when "001010001001" => q <= "00001011100010000000";
when "001010001010" => q <= "00001011100010000000";
when "001010001011" => q <= "00001011110010000000";
when "001010001100" => q <= "00001100000010000000";
when "001010001101" => q <= "00001100010010000000";
when "001010001110" => q <= "00001100110010000000";
when "001010001111" => q <= "00001101000010000000";
when "001010010000" => q <= "00001101100010000000";
when "001010010001" => q <= "00001101110010000000";
when "001010010010" => q <= "00001110010010000000";
when "001010010011" => q <= "00001110110010000000";
when "001010010100" => q <= "00001111010010000000";
when "001010010101" => q <= "00001111100010000000";
when "001010010110" => q <= "00010000000010000000";
when "001010010111" => q <= "00010000100010000000";
when "001010011000" => q <= "00010001000001111100";
when "001010011001" => q <= "00010001010001110111";
when "001010011010" => q <= "00010001110001110011";
when "001010011011" => q <= "00010010010001101110";
when "001010011100" => q <= "00010010110001101000";
when "001010011101" => q <= "00010011100001100010";
when "001010011110" => q <= "00010100000001011011";
when "001010011111" => q <= "00010100110001010011";
when "001010100000" => q <= "00010101100001001010";
when "001010100001" => q <= "00010110010001000000";
when "001010100010" => q <= "00010111000000110110";
when "001010100011" => q <= "00010111110000101011";
when "001010100100" => q <= "00011000100000100001";
when "001010100101" => q <= "00011000110000011011";
when "001010100110" => q <= "00011000110000011001";
when "001010100111" => q <= "00011000100000100000";
when "001011000000" => q <= "00000100000010000000";
when "001011000001" => q <= "00000101110010000000";
when "001011000010" => q <= "00000111010010000000";
when "001011000011" => q <= "00001000010010000000";
when "001011000100" => q <= "00001000110010000000";
when "001011000101" => q <= "00001001010010000000";
when "001011000110" => q <= "00001001100010000000";
when "001011000111" => q <= "00001001110010000000";
when "001011001000" => q <= "00001010000010000000";
when "001011001001" => q <= "00001010010010000000";
when "001011001010" => q <= "00001010100010000000";
when "001011001011" => q <= "00001010110010000000";
when "001011001100" => q <= "00001011000010000000";
when "001011001101" => q <= "00001011010010000000";
when "001011001110" => q <= "00001011110010000000";
when "001011001111" => q <= "00001100000010000000";
when "001011010000" => q <= "00001100100010000000";
when "001011010001" => q <= "00001101000010000000";
when "001011010010" => q <= "00001101010010000000";
when "001011010011" => q <= "00001101110010000000";
when "001011010100" => q <= "00001110010010000000";
when "001011010101" => q <= "00001110110010000000";
when "001011010110" => q <= "00001111000010000000";
when "001011010111" => q <= "00001111100001111110";
when "001011011000" => q <= "00010000000001111010";
when "001011011001" => q <= "00010000010001110110";
when "001011011010" => q <= "00010000110001110001";
when "001011011011" => q <= "00010001010001101100";
when "001011011100" => q <= "00010001110001100111";
when "001011011101" => q <= "00010010010001100001";
when "001011011110" => q <= "00010010110001011010";
when "001011011111" => q <= "00010011100001010010";
when "001011100000" => q <= "00010100000001001010";
when "001011100001" => q <= "00010100110001000000";
when "001011100010" => q <= "00010101100000110101";
when "001011100011" => q <= "00010110010000101010";
when "001011100100" => q <= "00010110110000100000";
when "001011100101" => q <= "00010111010000011000";
when "001011100110" => q <= "00010111100000010101";
when "001011100111" => q <= "00010111010000011011";
when "001100000000" => q <= "00000100000010000000";
when "001100000001" => q <= "00000101010010000000";
when "001100000010" => q <= "00000110010010000000";
when "001100000011" => q <= "00000111000010000000";
when "001100000100" => q <= "00000111100010000000";
when "001100000101" => q <= "00001000000010000000";
when "001100000110" => q <= "00001000010010000000";
when "001100000111" => q <= "00001000110010000000";
when "001100001000" => q <= "00001001000010000000";
when "001100001001" => q <= "00001001010010000000";
when "001100001010" => q <= "00001001100010000000";
when "001100001011" => q <= "00001001110010000000";
when "001100001100" => q <= "00001010000010000000";
when "001100001101" => q <= "00001010100010000000";
when "001100001110" => q <= "00001010110010000000";
when "001100001111" => q <= "00001011010010000000";
when "001100010000" => q <= "00001011100010000000";
when "001100010001" => q <= "00001100000010000000";
when "001100010010" => q <= "00001100100010000000";
when "001100010011" => q <= "00001101000010000000";
when "001100010100" => q <= "00001101010010000000";
when "001100010101" => q <= "00001101110010000000";
when "001100010110" => q <= "00001110000010000000";
when "001100010111" => q <= "00001110100001111101";
when "001100011000" => q <= "00001111000001111000";
when "001100011001" => q <= "00001111010001110100";
when "001100011010" => q <= "00001111110001110000";
when "001100011011" => q <= "00010000010001101011";
when "001100011100" => q <= "00010000110001100110";
when "001100011101" => q <= "00010001000001100000";
when "001100011110" => q <= "00010001110001011001";
when "001100011111" => q <= "00010010010001010001";
when "001100100000" => q <= "00010010110001001001";
when "001100100001" => q <= "00010011010000111111";
when "001100100010" => q <= "00010100000000110100";
when "001100100011" => q <= "00010100100000101001";
when "001100100100" => q <= "00010101000000011110";
when "001100100101" => q <= "00010101100000010110";
when "001100100110" => q <= "00010101110000010011";
when "001100100111" => q <= "00010101110000010111";
when "001101000000" => q <= "00000100000010000000";
when "001101000001" => q <= "00000100110010000000";
when "001101000010" => q <= "00000101100010000000";
when "001101000011" => q <= "00000110000010000000";
when "001101000100" => q <= "00000110010010000000";
when "001101000101" => q <= "00000110110010000000";
when "001101000110" => q <= "00000111010010000000";
when "001101000111" => q <= "00000111100010000000";
when "001101001000" => q <= "00000111110010000000";
when "001101001001" => q <= "00001000010010000000";
when "001101001010" => q <= "00001000100010000000";
when "001101001011" => q <= "00001000110010000000";
when "001101001100" => q <= "00001001010010000000";
when "001101001101" => q <= "00001001100010000000";
when "001101001110" => q <= "00001010000010000000";
when "001101001111" => q <= "00001010010010000000";
when "001101010000" => q <= "00001010110010000000";
when "001101010001" => q <= "00001011000010000000";
when "001101010010" => q <= "00001011100010000000";
when "001101010011" => q <= "00001100000010000000";
when "001101010100" => q <= "00001100010010000000";
when "001101010101" => q <= "00001100110010000000";
when "001101010110" => q <= "00001101010001111111";
when "001101010111" => q <= "00001101100001111011";
when "001101011000" => q <= "00001110000001110111";
when "001101011001" => q <= "00001110010001110010";
when "001101011010" => q <= "00001110110001101110";
when "001101011011" => q <= "00001111010001101001";
when "001101011100" => q <= "00001111100001100100";
when "001101011101" => q <= "00010000000001011110";
when "001101011110" => q <= "00010000100001011000";
when "001101011111" => q <= "00010001000001010000";
when "001101100000" => q <= "00010001100001000111";
when "001101100001" => q <= "00010010000000111101";
when "001101100010" => q <= "00010010100000110011";
when "001101100011" => q <= "00010011000000100111";
when "001101100100" => q <= "00010011100000011101";
when "001101100101" => q <= "00010011110000010100";
when "001101100110" => q <= "00010100010000010000";
when "001101100111" => q <= "00010100100000010011";
when "001110000000" => q <= "00000011110010000000";
when "001110000001" => q <= "00000100000010000000";
when "001110000010" => q <= "00000100010010000000";
when "001110000011" => q <= "00000100110010000000";
when "001110000100" => q <= "00000101000010000000";
when "001110000101" => q <= "00000101100010000000";
when "001110000110" => q <= "00000110000010000000";
when "001110000111" => q <= "00000110010010000000";
when "001110001000" => q <= "00000110110010000000";
when "001110001001" => q <= "00000111000010000000";
when "001110001010" => q <= "00000111100010000000";
when "001110001011" => q <= "00000111110010000000";
when "001110001100" => q <= "00001000010010000000";
when "001110001101" => q <= "00001000110010000000";
when "001110001110" => q <= "00001001000010000000";
when "001110001111" => q <= "00001001100010000000";
when "001110010000" => q <= "00001001110010000000";
when "001110010001" => q <= "00001010010010000000";
when "001110010010" => q <= "00001010100010000000";
when "001110010011" => q <= "00001011000010000000";
when "001110010100" => q <= "00001011010010000000";
when "001110010101" => q <= "00001011110010000000";
when "001110010110" => q <= "00001100010001111110";
when "001110010111" => q <= "00001100100001111001";
when "001110011000" => q <= "00001101000001110101";
when "001110011001" => q <= "00001101010001110001";
when "001110011010" => q <= "00001101110001101100";
when "001110011011" => q <= "00001110000001101000";
when "001110011100" => q <= "00001110100001100010";
when "001110011101" => q <= "00001110110001011101";
when "001110011110" => q <= "00001111010001010110";
when "001110011111" => q <= "00001111110001001111";
when "001110100000" => q <= "00010000000001000110";
when "001110100001" => q <= "00010000100000111100";
when "001110100010" => q <= "00010001000000110001";
when "001110100011" => q <= "00010001010000100110";
when "001110100100" => q <= "00010001110000011011";
when "001110100101" => q <= "00010010010000010010";
when "001110100110" => q <= "00010010100000001110";
when "001110100111" => q <= "00010011000000010001";
when "001111000000" => q <= "00000011100010000000";
when "001111000001" => q <= "00000011010010000000";
when "001111000010" => q <= "00000011010010000000";
when "001111000011" => q <= "00000011100010000000";
when "001111000100" => q <= "00000011110010000000";
when "001111000101" => q <= "00000100010010000000";
when "001111000110" => q <= "00000100110010000000";
when "001111000111" => q <= "00000101000010000000";
when "001111001000" => q <= "00000101100010000000";
when "001111001001" => q <= "00000110000010000000";
when "001111001010" => q <= "00000110100010000000";
when "001111001011" => q <= "00000111000010000000";
when "001111001100" => q <= "00000111010010000000";
when "001111001101" => q <= "00000111110010000000";
when "001111001110" => q <= "00001000000010000000";
when "001111001111" => q <= "00001000100010000000";
when "001111010000" => q <= "00001001000010000000";
when "001111010001" => q <= "00001001010010000000";
when "001111010010" => q <= "00001001100010000000";
when "001111010011" => q <= "00001010000010000000";
when "001111010100" => q <= "00001010010010000000";
when "001111010101" => q <= "00001010110010000000";
when "001111010110" => q <= "00001011000001111100";
when "001111010111" => q <= "00001011100001111000";
when "001111011000" => q <= "00001100000001110100";
when "001111011001" => q <= "00001100010001101111";
when "001111011010" => q <= "00001100110001101011";
when "001111011011" => q <= "00001101000001100110";
when "001111011100" => q <= "00001101100001100001";
when "001111011101" => q <= "00001101110001011011";
when "001111011110" => q <= "00001110000001010100";
when "001111011111" => q <= "00001110100001001101";
when "001111100000" => q <= "00001110110001000100";
when "001111100001" => q <= "00001111000000111010";
when "001111100010" => q <= "00001111100000101111";
when "001111100011" => q <= "00001111110000100100";
when "001111100100" => q <= "00010000000000011001";
when "001111100101" => q <= "00010000100000010001";
when "001111100110" => q <= "00010001000000001100";
when "001111100111" => q <= "00010001010000010000";
when "010000000000" => q <= "00000011010010000000";
when "010000000001" => q <= "00000010110010000000";
when "010000000010" => q <= "00000010010010000000";
when "010000000011" => q <= "00000010010010000000";
when "010000000100" => q <= "00000010100010000000";
when "010000000101" => q <= "00000011000010000000";
when "010000000110" => q <= "00000011100010000000";
when "010000000111" => q <= "00000100000010000000";
when "010000001000" => q <= "00000100100010000000";
when "010000001001" => q <= "00000101000010000000";
when "010000001010" => q <= "00000101100010000000";
when "010000001011" => q <= "00000110000010000000";
when "010000001100" => q <= "00000110100010000000";
when "010000001101" => q <= "00000110110010000000";
when "010000001110" => q <= "00000111010010000000";
when "010000001111" => q <= "00000111100010000000";
when "010000010000" => q <= "00001000000010000000";
when "010000010001" => q <= "00001000010010000000";
when "010000010010" => q <= "00001000110010000000";
when "010000010011" => q <= "00001001000010000000";
when "010000010100" => q <= "00001001010010000000";
when "010000010101" => q <= "00001001110001111111";
when "010000010110" => q <= "00001010000001111011";
when "010000010111" => q <= "00001010100001110110";
when "010000011000" => q <= "00001010110001110010";
when "010000011001" => q <= "00001011010001101110";
when "010000011010" => q <= "00001011100001101001";
when "010000011011" => q <= "00001100000001100100";
when "010000011100" => q <= "00001100010001011111";
when "010000011101" => q <= "00001100100001011001";
when "010000011110" => q <= "00001101000001010010";
when "010000011111" => q <= "00001101010001001011";
when "010000100000" => q <= "00001101100001000010";
when "010000100001" => q <= "00001101110000111000";
when "010000100010" => q <= "00001110000000101101";
when "010000100011" => q <= "00001110000000100010";
when "010000100100" => q <= "00001110100000010111";
when "010000100101" => q <= "00001110110000001111";
when "010000100110" => q <= "00001111010000001011";
when "010000100111" => q <= "00010000000000001111";
when "010001000000" => q <= "00000011010010000000";
when "010001000001" => q <= "00000010000010000000";
when "010001000010" => q <= "00000001100010000000";
when "010001000011" => q <= "00000001010010000000";
when "010001000100" => q <= "00000001010010000000";
when "010001000101" => q <= "00000001110010000000";
when "010001000110" => q <= "00000010010010000000";
when "010001000111" => q <= "00000010110010000000";
when "010001001000" => q <= "00000011010010000000";
when "010001001001" => q <= "00000011110010000000";
when "010001001010" => q <= "00000100100010000000";
when "010001001011" => q <= "00000101000010000000";
when "010001001100" => q <= "00000101100010000000";
when "010001001101" => q <= "00000101110010000000";
when "010001001110" => q <= "00000110010010000000";
when "010001001111" => q <= "00000110110010000000";
when "010001010000" => q <= "00000111000010000000";
when "010001010001" => q <= "00000111010010000000";
when "010001010010" => q <= "00000111110010000000";
when "010001010011" => q <= "00001000000010000000";
when "010001010100" => q <= "00001000100010000000";
when "010001010101" => q <= "00001000110001111101";
when "010001010110" => q <= "00001001000001111001";
when "010001010111" => q <= "00001001100001110101";
when "010001011000" => q <= "00001001110001110000";
when "010001011001" => q <= "00001010010001101100";
when "010001011010" => q <= "00001010100001100111";
when "010001011011" => q <= "00001010110001100010";
when "010001011100" => q <= "00001011010001011101";
when "010001011101" => q <= "00001011100001010111";
when "010001011110" => q <= "00001011110001010000";
when "010001011111" => q <= "00001011110001001000";
when "010001100000" => q <= "00001100000000111111";
when "010001100001" => q <= "00001100010000110101";
when "010001100010" => q <= "00001100010000101010";
when "010001100011" => q <= "00001100100000011111";
when "010001100100" => q <= "00001100110000010101";
when "010001100101" => q <= "00001101000000001101";
when "010001100110" => q <= "00001101100000001010";
when "010001100111" => q <= "00001110100000010000";
when "010010000000" => q <= "00000011110010000000";
when "010010000001" => q <= "00000001110010000000";
when "010010000010" => q <= "00000000110010000000";
when "010010000011" => q <= "00000000010010000000";
when "010010000100" => q <= "00000000000010000000";
when "010010000101" => q <= "00000000010010000000";
when "010010000110" => q <= "00000000110010000000";
when "010010000111" => q <= "00000001100010000000";
when "010010001000" => q <= "00000010000010000000";
when "010010001001" => q <= "00000010110010000000";
when "010010001010" => q <= "00000011010010000000";
when "010010001011" => q <= "00000011110010000000";
when "010010001100" => q <= "00000100100010000000";
when "010010001101" => q <= "00000101000010000000";
when "010010001110" => q <= "00000101010010000000";
when "010010001111" => q <= "00000101110010000000";
when "010010010000" => q <= "00000110000010000000";
when "010010010001" => q <= "00000110100010000000";
when "010010010010" => q <= "00000110110010000000";
when "010010010011" => q <= "00000111000010000000";
when "010010010100" => q <= "00000111100010000000";
when "010010010101" => q <= "00000111110001111100";
when "010010010110" => q <= "00001000000001110111";
when "010010010111" => q <= "00001000100001110011";
when "010010011000" => q <= "00001000110001101111";
when "010010011001" => q <= "00001001000001101010";
when "010010011010" => q <= "00001001100001100110";
when "010010011011" => q <= "00001001110001100001";
when "010010011100" => q <= "00001010000001011011";
when "010010011101" => q <= "00001010010001010101";
when "010010011110" => q <= "00001010010001001110";
when "010010011111" => q <= "00001010100001000110";
when "010010100000" => q <= "00001010100000111101";
when "010010100001" => q <= "00001010100000110011";
when "010010100010" => q <= "00001010110000101000";
when "010010100011" => q <= "00001010110000011101";
when "010010100100" => q <= "00001011000000010011";
when "010010100101" => q <= "00001011100000001100";
when "010010100110" => q <= "00001100000000001010";
when "010010100111" => q <= "00001101000000010001";
when "010011000000" => q <= "00000100100001110100";
when "010011000001" => q <= "00000001110010000000";
when "010011000010" => q <= "00000000000010000000";
when "010011000011" => q <= "00000000000010000000";
when "010011000100" => q <= "00000000000010000000";
when "010011000101" => q <= "00000000000010000000";
when "010011000110" => q <= "00000000000010000000";
when "010011000111" => q <= "00000000000010000000";
when "010011001000" => q <= "00000000110010000000";
when "010011001001" => q <= "00000001100010000000";
when "010011001010" => q <= "00000010000010000000";
when "010011001011" => q <= "00000010110010000000";
when "010011001100" => q <= "00000011010010000000";
when "010011001101" => q <= "00000011110010000000";
when "010011001110" => q <= "00000100010010000000";
when "010011001111" => q <= "00000100110010000000";
when "010011010000" => q <= "00000101000010000000";
when "010011010001" => q <= "00000101100010000000";
when "010011010010" => q <= "00000101110010000000";
when "010011010011" => q <= "00000110000010000000";
when "010011010100" => q <= "00000110100001111110";
when "010011010101" => q <= "00000110110001111010";
when "010011010110" => q <= "00000111000001110110";
when "010011010111" => q <= "00000111100001110010";
when "010011011000" => q <= "00000111110001101101";
when "010011011001" => q <= "00001000000001101001";
when "010011011010" => q <= "00001000010001100100";
when "010011011011" => q <= "00001000100001011111";
when "010011011100" => q <= "00001000110001011001";
when "010011011101" => q <= "00001001000001010010";
when "010011011110" => q <= "00001001000001001011";
when "010011011111" => q <= "00001001000001000011";
when "010011100000" => q <= "00001001000000111010";
when "010011100001" => q <= "00001001000000101111";
when "010011100010" => q <= "00001001000000100101";
when "010011100011" => q <= "00001001000000011010";
when "010011100100" => q <= "00001001010000010001";
when "010011100101" => q <= "00001001110000001011";
when "010011100110" => q <= "00001010100000001011";
when "010011100111" => q <= "00001100000000010100";
when "010100000000" => q <= "00000101110001100010";
when "010100000001" => q <= "00000010000010000000";
when "010100000010" => q <= "00000000000010000000";
when "010100000011" => q <= "00000000000010000000";
when "010100000100" => q <= "00000000000010000000";
when "010100000101" => q <= "00000000000010000000";
when "010100000110" => q <= "00000000000010000000";
when "010100000111" => q <= "00000000000010000000";
when "010100001000" => q <= "00000000000010000000";
when "010100001001" => q <= "00000000000010000000";
when "010100001010" => q <= "00000000110010000000";
when "010100001011" => q <= "00000001100010000000";
when "010100001100" => q <= "00000010000010000000";
when "010100001101" => q <= "00000010110010000000";
when "010100001110" => q <= "00000011010010000000";
when "010100001111" => q <= "00000011110010000000";
when "010100010000" => q <= "00000100000010000000";
when "010100010001" => q <= "00000100100010000000";
when "010100010010" => q <= "00000100110010000000";
when "010100010011" => q <= "00000101000010000000";
when "010100010100" => q <= "00000101100001111101";
when "010100010101" => q <= "00000101110001111001";
when "010100010110" => q <= "00000110000001110100";
when "010100010111" => q <= "00000110010001110000";
when "010100011000" => q <= "00000110110001101100";
when "010100011001" => q <= "00000111000001100111";
when "010100011010" => q <= "00000111010001100010";
when "010100011011" => q <= "00000111010001011100";
when "010100011100" => q <= "00000111100001010110";
when "010100011101" => q <= "00000111100001010000";
when "010100011110" => q <= "00000111100001001000";
when "010100011111" => q <= "00000111100001000000";
when "010100100000" => q <= "00000111100000110110";
when "010100100001" => q <= "00000111010000101100";
when "010100100010" => q <= "00000111010000100010";
when "010100100011" => q <= "00000111010000011000";
when "010100100100" => q <= "00000111100000001111";
when "010100100101" => q <= "00001000010000001011";
when "010100100110" => q <= "00001001010000001101";
when "010100100111" => q <= "00001011010000011010";
when "010101000000" => q <= "00000111110001001100";
when "010101000001" => q <= "00000011000010000000";
when "010101000010" => q <= "00000000000010000000";
when "010101000011" => q <= "00000000000010000000";
when "010101000100" => q <= "00000000000010000000";
when "010101000101" => q <= "00000000000010000000";
when "010101000110" => q <= "00000000000010000000";
when "010101000111" => q <= "00000000000010000000";
when "010101001000" => q <= "00000000000010000000";
when "010101001001" => q <= "00000000000010000000";
when "010101001010" => q <= "00000000000010000000";
when "010101001011" => q <= "00000000000010000000";
when "010101001100" => q <= "00000000110010000000";
when "010101001101" => q <= "00000001100010000000";
when "010101001110" => q <= "00000010000010000000";
when "010101001111" => q <= "00000010100010000000";
when "010101010000" => q <= "00000011000010000000";
when "010101010001" => q <= "00000011010010000000";
when "010101010010" => q <= "00000011110010000000";
when "010101010011" => q <= "00000100000001111111";
when "010101010100" => q <= "00000100010001111011";
when "010101010101" => q <= "00000100110001110111";
when "010101010110" => q <= "00000101000001110011";
when "010101010111" => q <= "00000101010001101110";
when "010101011000" => q <= "00000101100001101010";
when "010101011001" => q <= "00000101110001100101";
when "010101011010" => q <= "00000101110001100000";
when "010101011011" => q <= "00000110000001011010";
when "010101011100" => q <= "00000110000001010100";
when "010101011101" => q <= "00000110000001001101";
when "010101011110" => q <= "00000110000001000101";
when "010101011111" => q <= "00000101110000111100";
when "010101100000" => q <= "00000101110000110011";
when "010101100001" => q <= "00000101100000101001";
when "010101100010" => q <= "00000101100000011111";
when "010101100011" => q <= "00000101100000010101";
when "010101100100" => q <= "00000110000000001110";
when "010101100101" => q <= "00000110110000001100";
when "010101100110" => q <= "00001000010000010001";
when "010101100111" => q <= "00001010110000100001";
when "010110000000" => q <= "00001011000000110000";
when "010110000001" => q <= "00000100110001110011";
when "010110000010" => q <= "00000000100010000000";
when "010110000011" => q <= "00000000000010000000";
when "010110000100" => q <= "00000000000010000000";
when "010110000101" => q <= "00000000000010000000";
when "010110000110" => q <= "00000000000010000000";
when "010110000111" => q <= "00000000000010000000";
when "010110001000" => q <= "00000000000010000000";
when "010110001001" => q <= "00000000000010000000";
when "010110001010" => q <= "00000000000010000000";
when "010110001011" => q <= "00000000000010000000";
when "010110001100" => q <= "00000000000010000000";
when "010110001101" => q <= "00000000000010000000";
when "010110001110" => q <= "00000000110010000000";
when "010110001111" => q <= "00000001010010000000";
when "010110010000" => q <= "00000001110010000000";
when "010110010001" => q <= "00000010000010000000";
when "010110010010" => q <= "00000010100010000000";
when "010110010011" => q <= "00000010110001111110";
when "010110010100" => q <= "00000011010001111010";
when "010110010101" => q <= "00000011100001110101";
when "010110010110" => q <= "00000011110001110001";
when "010110010111" => q <= "00000100000001101101";
when "010110011000" => q <= "00000100010001101000";
when "010110011001" => q <= "00000100010001100011";
when "010110011010" => q <= "00000100100001011101";
when "010110011011" => q <= "00000100100001010111";
when "010110011100" => q <= "00000100100001010001";
when "010110011101" => q <= "00000100010001001010";
when "010110011110" => q <= "00000100010001000001";
when "010110011111" => q <= "00000100000000111001";
when "010110100000" => q <= "00000011110000101111";
when "010110100001" => q <= "00000011100000100101";
when "010110100010" => q <= "00000011100000011100";
when "010110100011" => q <= "00000011110000010011";
when "010110100100" => q <= "00000100100000001110";
when "010110100101" => q <= "00000101110000001110";
when "010110100110" => q <= "00000111110000010111";
when "010110100111" => q <= "00001010110000101100";
when "010111000000" => q <= "00001111100000001110";
when "010111000001" => q <= "00000111110001011010";
when "010111000010" => q <= "00000010000010000000";
when "010111000011" => q <= "00000000000010000000";
when "010111000100" => q <= "00000000000010000000";
when "010111000101" => q <= "00000000000010000000";
when "010111000110" => q <= "00000000000010000000";
when "010111000111" => q <= "00000000000010000000";
when "010111001000" => q <= "00000000000010000000";
when "010111001001" => q <= "00000000000010000000";
when "010111001010" => q <= "00000000000010000000";
when "010111001011" => q <= "00000000000010000000";
when "010111001100" => q <= "00000000000010000000";
when "010111001101" => q <= "00000000000010000000";
when "010111001110" => q <= "00000000000010000000";
when "010111001111" => q <= "00000000000010000000";
when "010111010000" => q <= "00000000010010000000";
when "010111010001" => q <= "00000000110010000000";
when "010111010010" => q <= "00000001010010000000";
when "010111010011" => q <= "00000001100001111101";
when "010111010100" => q <= "00000001110001111000";
when "010111010101" => q <= "00000010000001110100";
when "010111010110" => q <= "00000010010001101111";
when "010111010111" => q <= "00000010100001101011";
when "010111011000" => q <= "00000010110001100110";
when "010111011001" => q <= "00000010110001100000";
when "010111011010" => q <= "00000010110001011011";
when "010111011011" => q <= "00000010110001010100";
when "010111011100" => q <= "00000010110001001110";
when "010111011101" => q <= "00000010100001000110";
when "010111011110" => q <= "00000010010000111110";
when "010111011111" => q <= "00000010000000110101";
when "010111100000" => q <= "00000001110000101011";
when "010111100001" => q <= "00000001110000100010";
when "010111100010" => q <= "00000001110000011001";
when "010111100011" => q <= "00000010010000010011";
when "010111100100" => q <= "00000011010000010000";
when "010111100101" => q <= "00000101000000010011";
when "010111100110" => q <= "00000111110000100000";
when "010111100111" => q <= "00001011110000111100";
when "011000000000" => q <= "00010110000000000000";
when "011000000001" => q <= "00001100000000111010";
when "011000000010" => q <= "00000100110001110101";
when "011000000011" => q <= "00000000000010000000";
when "011000000100" => q <= "00000000000010000000";
when "011000000101" => q <= "00000000000010000000";
when "011000000110" => q <= "00000000000010000000";
when "011000000111" => q <= "00000000000010000000";
when "011000001000" => q <= "00000000000010000000";
when "011000001001" => q <= "00000000000010000000";
when "011000001010" => q <= "00000000000010000000";
when "011000001011" => q <= "00000000000010000000";
when "011000001100" => q <= "00000000000010000000";
when "011000001101" => q <= "00000000000010000000";
when "011000001110" => q <= "00000000000010000000";
when "011000001111" => q <= "00000000000010000000";
when "011000010000" => q <= "00000000000010000000";
when "011000010001" => q <= "00000000000010000000";
when "011000010010" => q <= "00000000000010000000";
when "011000010011" => q <= "00000000000001111011";
when "011000010100" => q <= "00000000010001110111";
when "011000010101" => q <= "00000000100001110010";
when "011000010110" => q <= "00000000110001101101";
when "011000010111" => q <= "00000001000001101001";
when "011000011000" => q <= "00000001000001100011";
when "011000011001" => q <= "00000001000001011110";
when "011000011010" => q <= "00000001000001011000";
when "011000011011" => q <= "00000001000001010001";
when "011000011100" => q <= "00000000110001001010";
when "011000011101" => q <= "00000000100001000010";
when "011000011110" => q <= "00000000010000111010";
when "011000011111" => q <= "00000000000000110001";
when "011000100000" => q <= "00000000000000101000";
when "011000100001" => q <= "00000000000000011111";
when "011000100010" => q <= "00000000010000011000";
when "011000100011" => q <= "00000001000000010011";
when "011000100100" => q <= "00000010100000010011";
when "011000100101" => q <= "00000100110000011011";
when "011000100110" => q <= "00001000100000101101";
when "011000100111" => q <= "00001110000001010000";
when "011001000000" => q <= "00011110110000000000";
when "011001000001" => q <= "00010010010000010010";
when "011001000010" => q <= "00001001000001010111";
when "011001000011" => q <= "00000010010010000000";
when "011001000100" => q <= "00000000000010000000";
when "011001000101" => q <= "00000000000010000000";
when "011001000110" => q <= "00000000000010000000";
when "011001000111" => q <= "00000000000010000000";
when "011001001000" => q <= "00000000000010000000";
when "011001001001" => q <= "00000000000010000000";
when "011001001010" => q <= "00000000000010000000";
when "011001001011" => q <= "00000000000010000000";
when "011001001100" => q <= "00000000000010000000";
when "011001001101" => q <= "00000000000010000000";
when "011001001110" => q <= "00000000000010000000";
when "011001001111" => q <= "00000000000010000000";
when "011001010000" => q <= "00000000000010000000";
when "011001010001" => q <= "00000000000010000000";
when "011001010010" => q <= "00000000000001111111";
when "011001010011" => q <= "00000000000001111010";
when "011001010100" => q <= "00000000000001110101";
when "011001010101" => q <= "00000000000001110001";
when "011001010110" => q <= "00000000000001101100";
when "011001010111" => q <= "00000000000001100110";
when "011001011000" => q <= "00000000000001100001";
when "011001011001" => q <= "00000000000001011011";
when "011001011010" => q <= "00000000000001010101";
when "011001011011" => q <= "00000000000001001110";
when "011001011100" => q <= "00000000000001000110";
when "011001011101" => q <= "00000000000000111111";
when "011001011110" => q <= "00000000000000110110";
when "011001011111" => q <= "00000000000000101101";
when "011001100000" => q <= "00000000000000100101";
when "011001100001" => q <= "00000000000000011101";
when "011001100010" => q <= "00000000000000011000";
when "011001100011" => q <= "00000000000000010110";
when "011001100100" => q <= "00000010010000011010";
when "011001100101" => q <= "00000101110000100110";
when "011001100110" => q <= "00001010110001000000";
when "011001100111" => q <= "00010001110001101100";
when "011010000000" => q <= "00100000000000000000";
when "011010000001" => q <= "00011011000000000000";
when "011010000010" => q <= "00001111010000110001";
when "011010000011" => q <= "00000110100001101001";
when "011010000100" => q <= "00000000100010000000";
when "011010000101" => q <= "00000000000010000000";
when "011010000110" => q <= "00000000000010000000";
when "011010000111" => q <= "00000000000010000000";
when "011010001000" => q <= "00000000000010000000";
when "011010001001" => q <= "00000000000010000000";
when "011010001010" => q <= "00000000000010000000";
when "011010001011" => q <= "00000000000010000000";
when "011010001100" => q <= "00000000000010000000";
when "011010001101" => q <= "00000000000010000000";
when "011010001110" => q <= "00000000000010000000";
when "011010001111" => q <= "00000000000010000000";
when "011010010000" => q <= "00000000000010000000";
when "011010010001" => q <= "00000000000010000000";
when "011010010010" => q <= "00000000000001111110";
when "011010010011" => q <= "00000000000001111001";
when "011010010100" => q <= "00000000000001110100";
when "011010010101" => q <= "00000000000001101111";
when "011010010110" => q <= "00000000000001101010";
when "011010010111" => q <= "00000000000001100100";
when "011010011000" => q <= "00000000000001011110";
when "011010011001" => q <= "00000000000001011000";
when "011010011010" => q <= "00000000000001010001";
when "011010011011" => q <= "00000000000001001010";
when "011010011100" => q <= "00000000000001000011";
when "011010011101" => q <= "00000000000000111011";
when "011010011110" => q <= "00000000000000110011";
when "011010011111" => q <= "00000000000000101011";
when "011010100000" => q <= "00000000000000100011";
when "011010100001" => q <= "00000000000000011101";
when "011010100010" => q <= "00000000000000011010";
when "011010100011" => q <= "00000000000000011100";
when "011010100100" => q <= "00000011000000100100";
when "011010100101" => q <= "00000111110000110111";
when "011010100110" => q <= "00001110100001011001";
when "011010100111" => q <= "00010111100010000000";
when "011011000000" => q <= "00100000000000000000";
when "011011000001" => q <= "00100000000000000000";
when "011011000010" => q <= "00011000010000000010";
when "011011000011" => q <= "00001101000001000110";
when "011011000100" => q <= "00000100110001110100";
when "011011000101" => q <= "00000000000010000000";
when "011011000110" => q <= "00000000000010000000";
when "011011000111" => q <= "00000000000010000000";
when "011011001000" => q <= "00000000000010000000";
when "011011001001" => q <= "00000000000010000000";
when "011011001010" => q <= "00000000000010000000";
when "011011001011" => q <= "00000000000010000000";
when "011011001100" => q <= "00000000000010000000";
when "011011001101" => q <= "00000000000010000000";
when "011011001110" => q <= "00000000000010000000";
when "011011001111" => q <= "00000000000010000000";
when "011011010000" => q <= "00000000000010000000";
when "011011010001" => q <= "00000000000010000000";
when "011011010010" => q <= "00000000000001111101";
when "011011010011" => q <= "00000000000001111000";
when "011011010100" => q <= "00000000000001110011";
when "011011010101" => q <= "00000000000001101101";
when "011011010110" => q <= "00000000000001100111";
when "011011010111" => q <= "00000000000001100010";
when "011011011000" => q <= "00000000000001011100";
when "011011011001" => q <= "00000000000001010101";
when "011011011010" => q <= "00000000000001001110";
when "011011011011" => q <= "00000000000001000111";
when "011011011100" => q <= "00000000000000111111";
when "011011011101" => q <= "00000000000000111000";
when "011011011110" => q <= "00000000000000110000";
when "011011011111" => q <= "00000000000000101001";
when "011011100000" => q <= "00000000000000100011";
when "011011100001" => q <= "00000000000000011111";
when "011011100010" => q <= "00000000000000011111";
when "011011100011" => q <= "00000001000000100101";
when "011011100100" => q <= "00000101100000110100";
when "011011100101" => q <= "00001011110001001111";
when "011011100110" => q <= "00010100100001111011";
when "011011100111" => q <= "00100000000010000000";
when "011100000000" => q <= "00100000000000000000";
when "011100000001" => q <= "00100000000000000000";
when "011100000010" => q <= "00100000000000000000";
when "011100000011" => q <= "00010110110000011000";
when "011100000100" => q <= "00001011110001010010";
when "011100000101" => q <= "00000011110001111000";
when "011100000110" => q <= "00000000000010000000";
when "011100000111" => q <= "00000000000010000000";
when "011100001000" => q <= "00000000000010000000";
when "011100001001" => q <= "00000000000010000000";
when "011100001010" => q <= "00000000000010000000";
when "011100001011" => q <= "00000000000010000000";
when "011100001100" => q <= "00000000000010000000";
when "011100001101" => q <= "00000000000010000000";
when "011100001110" => q <= "00000000000010000000";
when "011100001111" => q <= "00000000000010000000";
when "011100010000" => q <= "00000000000010000000";
when "011100010001" => q <= "00000000000010000000";
when "011100010010" => q <= "00000000000001111101";
when "011100010011" => q <= "00000000000001110111";
when "011100010100" => q <= "00000000000001110001";
when "011100010101" => q <= "00000000000001101011";
when "011100010110" => q <= "00000000000001100101";
when "011100010111" => q <= "00000000000001011111";
when "011100011000" => q <= "00000000000001011001";
when "011100011001" => q <= "00000000000001010010";
when "011100011010" => q <= "00000000000001001011";
when "011100011011" => q <= "00000000000001000100";
when "011100011100" => q <= "00000000000000111101";
when "011100011101" => q <= "00000000000000110101";
when "011100011110" => q <= "00000000000000101111";
when "011100011111" => q <= "00000000000000101001";
when "011100100000" => q <= "00000000000000100101";
when "011100100001" => q <= "00000000000000100101";
when "011100100010" => q <= "00000000000000101001";
when "011100100011" => q <= "00000011110000110101";
when "011100100100" => q <= "00001010000001001011";
when "011100100101" => q <= "00010010010001101111";
when "011100100110" => q <= "00011101110010000000";
when "011100100111" => q <= "00100000000010000000";
when "011101000000" => q <= "00100000000000000000";
when "011101000001" => q <= "00100000000000000000";
when "011101000010" => q <= "00100000000000000000";
when "011101000011" => q <= "00100000000000000000";
when "011101000100" => q <= "00010110000000100101";
when "011101000101" => q <= "00001011100001010111";
when "011101000110" => q <= "00000011100001111000";
when "011101000111" => q <= "00000000000010000000";
when "011101001000" => q <= "00000000000010000000";
when "011101001001" => q <= "00000000000010000000";
when "011101001010" => q <= "00000000000010000000";
when "011101001011" => q <= "00000000000010000000";
when "011101001100" => q <= "00000000000010000000";
when "011101001101" => q <= "00000000000010000000";
when "011101001110" => q <= "00000000000010000000";
when "011101001111" => q <= "00000000000010000000";
when "011101010000" => q <= "00000000000010000000";
when "011101010001" => q <= "00000000000010000000";
when "011101010010" => q <= "00000000000001111100";
when "011101010011" => q <= "00000000000001110110";
when "011101010100" => q <= "00000000000001110000";
when "011101010101" => q <= "00000000000001101010";
when "011101010110" => q <= "00000000000001100011";
when "011101010111" => q <= "00000000000001011101";
when "011101011000" => q <= "00000000000001010110";
when "011101011001" => q <= "00000000000001010000";
when "011101011010" => q <= "00000000000001001001";
when "011101011011" => q <= "00000000000001000010";
when "011101011100" => q <= "00000000000000111011";
when "011101011101" => q <= "00000000000000110101";
when "011101011110" => q <= "00000000000000101111";
when "011101011111" => q <= "00000000000000101100";
when "011101100000" => q <= "00000000000000101011";
when "011101100001" => q <= "00000000000000101110";
when "011101100010" => q <= "00000010110000111000";
when "011101100011" => q <= "00001000110001001011";
when "011101100100" => q <= "00010001010001101010";
when "011101100101" => q <= "00011100010010000000";
when "011101100110" => q <= "00100000000010000000";
when "011101100111" => q <= "00100000000010000000";

      when others => q <=   "00000000000000000000";
    end case;
  end process;

end rtl;

