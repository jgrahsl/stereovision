library ieee;
use ieee.std_logic_1164.all;
use IEEE.NUMERIC_STD.all;

library work;
use work.cam_pkg.all;

entity null_filter is
  generic (
    ID : integer range 0 to 63 := 0);
  port (
    pipe_in  : in  pipe_t;
    pipe_out : out pipe_t);
end null_filter;

architecture impl of null_filter is

  signal clk        : std_logic;
  signal rst        : std_logic;
  signal stage      : stage_t;
  signal stage_next : stage_t;

begin
  clk <= pipe_in.ctrl.clk;
  rst <= pipe_in.ctrl.rst;

  pipe_out.ctrl  <= pipe_in.ctrl;
  pipe_out.cfg   <= pipe_in.cfg;
  pipe_out.stage <= stage;

  process (pipe_in)
  begin
    stage_next <= pipe_in.stage;
  end process;

  proc_clk : process(pipe_in)
  begin
    if rst = '1' then
      stage.valid <= '0';
      stage.init  <= '0';
    else
      if rising_edge(clk) then
        if (pipe_in.cfg(ID).enable = '1') then
          stage <= stage_next;
        else
          stage <= pipe_in.stage;
        end if;
      end if;
    end if;
  end process;

end impl;
