../sim_pkg_32x32.vhd